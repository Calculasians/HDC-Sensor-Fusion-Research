`ifndef CONST
`define CONST

`define HV_DIMENSION 2000
`define CHANNEL_WIDTH 2
`define NGRAM_SIZE 3
`define TOTAL_NUM_CHANNEL 214
`define GSR_SRAM_ADDR_WIDTH 5
`define ECG_SRAM_ADDR_WIDTH 7
`define EEG_SRAM_ADDR_WIDTH 7
`define GSR_NUM_CHANNEL 32
`define ECG_NUM_CHANNEL 77
`define EEG_NUM_CHANNEL 105

`define ceilLog2(x) ( \
(x) > 2**30 ? 31 : \
(x) > 2**29 ? 30 : \
(x) > 2**28 ? 29 : \
(x) > 2**27 ? 28 : \
(x) > 2**26 ? 27 : \
(x) > 2**25 ? 26 : \
(x) > 2**24 ? 25 : \
(x) > 2**23 ? 24 : \
(x) > 2**22 ? 23 : \
(x) > 2**21 ? 22 : \
(x) > 2**20 ? 21 : \
(x) > 2**19 ? 20 : \
(x) > 2**18 ? 19 : \
(x) > 2**17 ? 18 : \
(x) > 2**16 ? 17 : \
(x) > 2**15 ? 16 : \
(x) > 2**14 ? 15 : \
(x) > 2**13 ? 14 : \
(x) > 2**12 ? 13 : \
(x) > 2**11 ? 12 : \
(x) > 2**10 ? 11 : \
(x) > 2**9 ? 10 : \
(x) > 2**8 ? 9 : \
(x) > 2**7 ? 8 : \
(x) > 2**6 ? 7 : \
(x) > 2**5 ? 6 : \
(x) > 2**4 ? 5 : \
(x) > 2**3 ? 4 : \
(x) > 2**2 ? 3 : \
(x) > 2**1 ? 2 : \
(x) > 2**0 ? 1 : 0)

`define IM_CHANNEL_TO_INDEX(i) ( \
(i) == 0 ? 16 : \
(i) == 1 ? 1 : \
(i) == 2 ? 8 : \
(i) == 3 ? 10 : \
(i) == 4 ? 3 : \
(i) == 5 ? 18 : \
(i) == 6 ? 12 : \
(i) == 7 ? 5 : \
(i) == 8 ? 20 : \
(i) == 9 ? 14 : \
(i) == 10 ? 0 : \
(i) == 11 ? 9 : \
(i) == 12 ? 2 : \
(i) == 13 ? 17 : \
(i) == 14 ? 11 : \
(i) == 15 ? 4 : \
(i) == 16 ? 19 : \
(i) == 17 ? 13 : \
(i) == 18 ? 6 : \
(i) == 19 ? 21 : \
(i) == 20 ? 1 : \
(i) == 21 ? 8 : \
(i) == 22 ? 16 : \
(i) == 23 ? 10 : \
(i) == 24 ? 3 : \
(i) == 25 ? 18 : \
(i) == 26 ? 12 : \
(i) == 27 ? 5 : \
(i) == 28 ? 20 : \
(i) == 29 ? 9 : \
(i) == 30 ? 0 : \
(i) == 31 ? 2 : \
(i) == 32 ? 17 : \
(i) == 33 ? 11 : \
(i) == 34 ? 4 : \
(i) == 35 ? 19 : \
(i) == 36 ? 13 : \
(i) == 37 ? 6 : \
(i) == 38 ? 8 : \
(i) == 39 ? 1 : \
(i) == 40 ? 16 : \
(i) == 41 ? 10 : \
(i) == 42 ? 3 : \
(i) == 43 ? 18 : \
(i) == 44 ? 12 : \
(i) == 45 ? 5 : \
(i) == 46 ? 17 : \
(i) == 47 ? 9 : \
(i) == 48 ? 2 : \
(i) == 49 ? 0 : \
(i) == 50 ? 11 : \
(i) == 51 ? 4 : \
(i) == 52 ? 19 : \
(i) == 53 ? 13 : \
(i) == 54 ? 16 : \
(i) == 55 ? 1 : \
(i) == 56 ? 8 : \
(i) == 57 ? 10 : \
(i) == 58 ? 3 : \
(i) == 59 ? 18 : \
(i) == 60 ? 12 : \
(i) == 61 ? 0 : \
(i) == 62 ? 9 : \
(i) == 63 ? 2 : \
(i) == 64 ? 17 : \
(i) == 65 ? 11 : \
(i) == 66 ? 4 : \
(i) == 67 ? 19 : \
(i) == 68 ? 1 : \
(i) == 69 ? 8 : \
(i) == 70 ? 16 : \
(i) == 71 ? 10 : \
(i) == 72 ? 3 : \
(i) == 73 ? 18 : \
(i) == 74 ? 9 : \
(i) == 75 ? 0 : \
(i) == 76 ? 2 : \
(i) == 77 ? 17 : \
(i) == 78 ? 11 : \
(i) == 79 ? 4 : \
(i) == 80 ? 8 : \
(i) == 81 ? 1 : \
(i) == 82 ? 16 : \
(i) == 83 ? 10 : \
(i) == 84 ? 3 : \
(i) == 85 ? 17 : \
(i) == 86 ? 9 : \
(i) == 87 ? 2 : \
(i) == 88 ? 0 : \
(i) == 89 ? 11 : \
(i) == 90 ? 16 : \
(i) == 91 ? 1 : \
(i) == 92 ? 8 : \
(i) == 93 ? 10 : \
(i) == 94 ? 0 : \
(i) == 95 ? 9 : \
(i) == 96 ? 2 : \
(i) == 97 ? 17 : \
(i) == 98 ? 1 : \
(i) == 99 ? 8 : \
(i) == 100 ? 16 : \
(i) == 101 ? 9 : \
(i) == 102 ? 0 : \
(i) == 103 ? 2 : \
(i) == 104 ? 8 : 0)

`define PROJM_POS_CHANNEL_TO_INDEX(i) ( \
(i) < 10 ? 15 : \
(i) < 20 ? 22 : \
(i) < 29 ? 21 : \
(i) < 38 ? 7 : \
(i) < 46 ? 6 : \
(i) < 54 ? 14 : \
(i) < 61 ? 13 : \
(i) < 68 ? 20 : \
(i) < 74 ? 19 : \
(i) < 80 ? 5 : \
(i) < 85 ? 4 : \
(i) < 90 ? 12 : \
(i) < 94 ? 11 : \
(i) < 98 ? 18 : \
(i) < 101 ? 17 : \
(i) < 104 ? 3 : \
(i) < 106 ? 2 : 0)

`define PROJM_NEG_CHANNEL_TO_INDEX(i) ( \
(i) < 10 ? 7 : \
(i) < 20 ? 15 : \
(i) < 29 ? 14 : \
(i) < 38 ? 21 : \
(i) < 46 ? 20 : \
(i) < 54 ? 6 : \
(i) < 61 ? 5 : \
(i) < 68 ? 13 : \
(i) < 74 ? 12 : \
(i) < 80 ? 19 : \
(i) < 85 ? 18 : \
(i) < 90 ? 4 : \
(i) < 94 ? 3 : \
(i) < 98 ? 11 : \
(i) < 101 ? 10 : \
(i) < 104 ? 17 : \
(i) < 106 ? 16 : 0)

`define PROTOTYPE_V_PLUS 2000'b01010111000011111010010011001101001110110101000000110001000000011011011101000100100110011000111111100100001010000100001010100011110000101110111111100011011100011011110010001001010001010111111011010001100011100111001101110100100001001001101001101011011001000000000010001110110010001010011101101001000110010100001100000010001100011101000100100011111110101110101101010010011110011100001111011000011101010000101111010101011111011011100100001111111001100110101101010101011101010001111100111001100011100011100101111000111111000111101101000101110111111110000010001010001111100000111101111010110000000101110101001100111110000110100110010000011111001111011100101011000110001011101101110100000100011000101101001111000001001111100101010000110010001101100111011010110000100001001111011000011001000010011000110001011010111110000001110110100000010011000100101001100101000100100101101001011011011101001010100111111010001110110101010111010110111011100100001010100011110011001101110010111111111010010110001001111000111110000000010011001010100111001011111111001100111000010101001100000001011100110110100000111001101001000100100010011011011111000001110100011011101101111101011011010100100110010000100000101110110101000110100001101111010111110011110101001010100100110100001111010001000100001100011011010110010100100101011100010100100000111001010000100101100001110110101100010001110101011000111001100010010100010111101000111110110001001001000011000100100000110011111000011110101001111010101110101111001100001000100111111010101111110010010010110010001101010111001001001100001111000000100011010010101110011100000110000100010011111010001110100110101001110011000100101101100110001110000011111101111000110010010011011100101100111110100100011110010110101101100000001101101101100110101100010011110001001111000000111000011001001000111000001111001100011101010100110001011010111100011101001010100111111101000011111111000010000101011110100011101011111111011010000100000110000011011100010110100110101100011101111001100101110010010001

`define PROTOTYPE_V_MIN 2000'b01010111000011111010000011001101001110111110000000110001000000011011011101000100101001111001011111100100001010000100000110100011000001001110111111011011000111011011110010001001010000010111111011010001110100000111001010110100100001001001100110101011011001000000000001001010110010001000011101110101000010010101111100000010001100011101000100000011111110101110101101010010011110011100001000011000101100000000101111000001011111011011100100000001001001100110101101010101011101010001111100111001100010001111010010011000111111100111101100110101110111111110000010001010000001111100111101111010110111000101111101001110110000000111100110000001111111001111011100101001000110001011101101100100110100000000101101111111000001001111011101010000111011101101100110101010110000100001001111011000010001000010011000110001001010010101011001110111100000010011000100101001010101100110101011100001011010111101111010101001111010001110110111010110110110110011100001010110100011110011000001110011000011111001110110001001111000111110000010010011001010100111001010011111001100111000010101001100011100111100110110100100111010001101000100100010010011010001000010110100011011101101111101011011010111010110010000100000101101001101000110100001101111101111110011110101101010100100110101111111010010000100001111111011010110010100100101100100010100100110111001010000101010110101110110101100010001100101011000111001100010010100010111001000111100110001001001000011000100100000110000101010011001111001111011001110101111001011001000100111111100101111110010010000110010001101010111001000001100001111000000100011010010110110001100000110000100010011011010001110100110101001110010111010101101100101101110001011111101111000110010010100011100101100111110100100011110010110101101100000010111100101100110101100010011110001001000101100100110011001001000110000000011001100011101010100110001011001111100101101001010010111111101000011111111111010100001011110100011101011000111011001100101000110000011011100010110100100101100011101111100000101110010101001

`define PROTOTYPE_A_HIGH 2000'b01010111000011111010010110001101001110110110000000110001000000011011011101000101100111110001011111100100001010000100000010110111110011001110111111011011011100011011111110001001010000010111111011010001101100000111001100110100100001001001111001101011011001000000000010101110110010001000011101110101000010001100001100000010001100011101000100100011111110101110101101010010011110011100001001011000100111010000101100101001011111011011010100000001111001100110101101010101011101010001111100111001100011101111010101011000111111100111101100100101110111111110000010001010001001100100111101111010110000010101111001001111110000000111100110010001111111001111011100101001000110001011101100010100001100000000101101110111000001001111011101010000111010011101100111011010110000100001001111011000011001000010011000110001001110000101001001110111101000010011000100101001010101101110101011101001011010111101111010100111111010000010110111010100110110111011100001010110100011110011101001110011000011111010010110001001111000111110000010010011001010100111001010011111001100111000010101001100000001111100110110100000111011010101000100100010010011011111000010110110011011101101111101011011010111000110010000100000101101001101000110100001101111101111110011110101001010100101110100001111010000000100001111111011010110010100100101011100000100100010111001010000101010100101110110101100010001100101011000111001100010010100010111011000110110110001001001000011000100100000110100111100011111111000111001001110101111001100001000100111111110101111110010010010110010010101010111001010001100001111000000100011010010110110011100110110000100010011011010001010100110101001110011000100101101100100101110000010111101111000110010010011011100101100111110100100011110010110101101100111001100000101100110101100010011110001001110101000100100011001001000111010010011001100011101010100110001011010111100101101001010010111111101000011111011000011110000011110100011101011111111011001100100100110000011011100010110100100101100011101111000010101110010101001

`define PROTOTYPE_A_LOW 2000'b01010111000011111010010101001101001110110101000000110001000000011011011101000100101110011001011111100100001010000100001110100011110000101110111111100011011110011011110010001001010011010111111011010001110111100111001010110100100101001001100010101011011001000000000010001110110010001011011101101001000000010010001100000010001100011101000101010011111110101110101101010010011110011100000001011000101111010000101111010101011111011011100100000001111001100110101001010101011101101001111100111001100011100011100000111000111111000111101101000001110111111110000010001010000001110000111101111010110111000101111101001110111110000111100110010011011100101111011100101001000110001011101101100100110100011000101101000111000001001111100101010000111010101101100111011010110000100001001011011000011001000010011000110001011010111110011101110111100000010011000100101001110101011110100011101001011011011100111010100111111010011110110101010101010110110011100000000010011011110011010001110011001110011001110100001001111000111110000001010011001010100111001011011111001100111000010101001100111010011100110110100100111000110111000100100010011111011111000010110100011011101101111101011011010110100110010000100000101001101101000110100001101111101111110011110101001010100100110100111111010011100100001100011011010101110100100101011100010100100110111001010000101001110100010110101100010001100101011000111001100010010100010111101000111000110001001001000011000100100000110011101010011000111001111010101110101111001001001011100111110010101111110010010101110010111101010111001101001100001111000000100011010010001111101100000110110100010011011010001100100110101001110001111010101101100110111110001011111101111000110010010011011100101100111110100100010110010110101101100000001101100101100110101100010011110000111100101000111000011001001000110100001111001111111101010100110001011001111100101101001010000111111101000011111111111010000111011110100011101011100111011001100101000110000011011100010110100010101100011101111001100101110010010001

`endif

