`ifndef CONST
`define CONST

`define HV_DIMENSION 2000
`define CHANNEL_WIDTH 2
`define NGRAM_SIZE 3
`define TOTAL_NUM_CHANNEL 214
`define GSR_SRAM_ADDR_WIDTH 5
`define ECG_SRAM_ADDR_WIDTH 7
`define EEG_SRAM_ADDR_WIDTH 7
`define GSR_NUM_CHANNEL 32
`define ECG_NUM_CHANNEL 77
`define EEG_NUM_CHANNEL 105

`define ceilLog2(x) ( \
(x) > 2**30 ? 31 : \
(x) > 2**29 ? 30 : \
(x) > 2**28 ? 29 : \
(x) > 2**27 ? 28 : \
(x) > 2**26 ? 27 : \
(x) > 2**25 ? 26 : \
(x) > 2**24 ? 25 : \
(x) > 2**23 ? 24 : \
(x) > 2**22 ? 23 : \
(x) > 2**21 ? 22 : \
(x) > 2**20 ? 21 : \
(x) > 2**19 ? 20 : \
(x) > 2**18 ? 19 : \
(x) > 2**17 ? 18 : \
(x) > 2**16 ? 17 : \
(x) > 2**15 ? 16 : \
(x) > 2**14 ? 15 : \
(x) > 2**13 ? 14 : \
(x) > 2**12 ? 13 : \
(x) > 2**11 ? 12 : \
(x) > 2**10 ? 11 : \
(x) > 2**9 ? 10 : \
(x) > 2**8 ? 9 : \
(x) > 2**7 ? 8 : \
(x) > 2**6 ? 7 : \
(x) > 2**5 ? 6 : \
(x) > 2**4 ? 5 : \
(x) > 2**3 ? 4 : \
(x) > 2**2 ? 3 : \
(x) > 2**1 ? 2 : \
(x) > 2**0 ? 1 : 0)

`define IM_CHANNEL_TO_INDEX(i) ( \
(i) == 0 ? 16 : \
(i) == 1 ? 1 : \
(i) == 2 ? 8 : \
(i) == 3 ? 10 : \
(i) == 4 ? 3 : \
(i) == 5 ? 18 : \
(i) == 6 ? 12 : \
(i) == 7 ? 5 : \
(i) == 8 ? 20 : \
(i) == 9 ? 14 : \
(i) == 10 ? 0 : \
(i) == 11 ? 9 : \
(i) == 12 ? 2 : \
(i) == 13 ? 17 : \
(i) == 14 ? 11 : \
(i) == 15 ? 4 : \
(i) == 16 ? 19 : \
(i) == 17 ? 13 : \
(i) == 18 ? 6 : \
(i) == 19 ? 21 : \
(i) == 20 ? 1 : \
(i) == 21 ? 8 : \
(i) == 22 ? 16 : \
(i) == 23 ? 10 : \
(i) == 24 ? 3 : \
(i) == 25 ? 18 : \
(i) == 26 ? 12 : \
(i) == 27 ? 5 : \
(i) == 28 ? 20 : \
(i) == 29 ? 9 : \
(i) == 30 ? 0 : \
(i) == 31 ? 2 : \
(i) == 32 ? 17 : \
(i) == 33 ? 11 : \
(i) == 34 ? 4 : \
(i) == 35 ? 19 : \
(i) == 36 ? 13 : \
(i) == 37 ? 6 : \
(i) == 38 ? 8 : \
(i) == 39 ? 1 : \
(i) == 40 ? 16 : \
(i) == 41 ? 10 : \
(i) == 42 ? 3 : \
(i) == 43 ? 18 : \
(i) == 44 ? 12 : \
(i) == 45 ? 5 : \
(i) == 46 ? 17 : \
(i) == 47 ? 9 : \
(i) == 48 ? 2 : \
(i) == 49 ? 0 : \
(i) == 50 ? 11 : \
(i) == 51 ? 4 : \
(i) == 52 ? 19 : \
(i) == 53 ? 13 : \
(i) == 54 ? 16 : \
(i) == 55 ? 1 : \
(i) == 56 ? 8 : \
(i) == 57 ? 10 : \
(i) == 58 ? 3 : \
(i) == 59 ? 18 : \
(i) == 60 ? 12 : \
(i) == 61 ? 0 : \
(i) == 62 ? 9 : \
(i) == 63 ? 2 : \
(i) == 64 ? 17 : \
(i) == 65 ? 11 : \
(i) == 66 ? 4 : \
(i) == 67 ? 19 : \
(i) == 68 ? 1 : \
(i) == 69 ? 8 : \
(i) == 70 ? 16 : \
(i) == 71 ? 10 : \
(i) == 72 ? 3 : \
(i) == 73 ? 18 : \
(i) == 74 ? 9 : \
(i) == 75 ? 0 : \
(i) == 76 ? 2 : \
(i) == 77 ? 17 : \
(i) == 78 ? 11 : \
(i) == 79 ? 4 : \
(i) == 80 ? 8 : \
(i) == 81 ? 1 : \
(i) == 82 ? 16 : \
(i) == 83 ? 10 : \
(i) == 84 ? 3 : \
(i) == 85 ? 17 : \
(i) == 86 ? 9 : \
(i) == 87 ? 2 : \
(i) == 88 ? 0 : \
(i) == 89 ? 11 : \
(i) == 90 ? 16 : \
(i) == 91 ? 1 : \
(i) == 92 ? 8 : \
(i) == 93 ? 10 : \
(i) == 94 ? 0 : \
(i) == 95 ? 9 : \
(i) == 96 ? 2 : \
(i) == 97 ? 17 : \
(i) == 98 ? 1 : \
(i) == 99 ? 8 : \
(i) == 100 ? 16 : \
(i) == 101 ? 9 : \
(i) == 102 ? 0 : \
(i) == 103 ? 2 : \
(i) == 104 ? 8 : 0)

`define PROJM_POS_CHANNEL_TO_INDEX(i) ( \
(i) < 10 ? 15 : \
(i) < 20 ? 22 : \
(i) < 29 ? 21 : \
(i) < 38 ? 7 : \
(i) < 46 ? 6 : \
(i) < 54 ? 14 : \
(i) < 61 ? 13 : \
(i) < 68 ? 20 : \
(i) < 74 ? 19 : \
(i) < 80 ? 5 : \
(i) < 85 ? 4 : \
(i) < 90 ? 12 : \
(i) < 94 ? 11 : \
(i) < 98 ? 18 : \
(i) < 101 ? 17 : \
(i) < 104 ? 3 : \
(i) < 106 ? 2 : 0)

`define PROJM_NEG_CHANNEL_TO_INDEX(i) ( \
(i) < 10 ? 7 : \
(i) < 20 ? 15 : \
(i) < 29 ? 14 : \
(i) < 38 ? 21 : \
(i) < 46 ? 20 : \
(i) < 54 ? 6 : \
(i) < 61 ? 5 : \
(i) < 68 ? 13 : \
(i) < 74 ? 12 : \
(i) < 80 ? 19 : \
(i) < 85 ? 18 : \
(i) < 90 ? 4 : \
(i) < 94 ? 3 : \
(i) < 98 ? 11 : \
(i) < 101 ? 10 : \
(i) < 104 ? 17 : \
(i) < 106 ? 16 : 0)

`define PROTOTYPE_V_PLUS 2000'b00111011010010110000110101010010010100111110111001110100011000101111000111101010100111101010010010001111110001011110100001100100010100010111111100100100010100011101011100000000111011011011010101001010000100111100011110110000000101110100010010000111001101110011011100110000101101001101010011111011110100110101000001110111011100110001110001111000101100111111001111011001010111010011111010100000010110110010111010001000001100000100111011010111110001100110010101011110101100001111101011110011100011100100001101111000111111101100000001101110010111011110001110001001100100111001000101011101110010110111110010100001011011101101101010100101000100110001010000101011111111101010011010101011100001111000010100011010111110000101010000000100010101110110100011011010011001001000100011011111000110111001001100100001111000110111011110011010011100111000111110000001010001110001000110011000011011111100000010001110110010101011010101000000101010001011101001100110000010010111100010000111110101010001011000010101001111001110100000100101100101100010011010001111001001100101010100000110101101100010000111110100000011101100000011100101101100010101100101001101100001101000010010011011010001010011000100100110010100000111100100101111001000001011011001101010010001011011110111001101001010001000000111111110110100011011001001111010101110010101101000011100011110111111010010101101001111001101101001100011101101011001110011010101111011100101010111011001011101001000101101110001111011001010111001010110010000111001111001010000011011010111110000000001101101001100001010100100000001100011001100101001001011000100000010100011000010111111010001100111111000110100001000011010000100101010011001101000011010110000001001010101001111100000111001000001110000000000110111011011011100101100001000000000001000001100001011001100010111111011011100011010101011101010110101111110110000101000000000000111010000010100100111100000101100000000110101010110010101010110110000011011111110110110110010000101010010100110000101011010010111101111101000000000

`define PROTOTYPE_V_MIN 2000'b00111011010001110000110100100010010100011110111000010100011000101111000111101010100111101010010010001111110001011111100001100100010101100111111100000100010101111101011100000000000011011011010101001010000100010100011110110000000101110100010010000111001111110011011100110000110101001101010011111011010100110110100001110111011100110001001011111000101100111111001111011001010001010011111010100000010001110010111010001000001101000110111011010111110001100110010101011110101101001111101011101111100011100100001101111000111111101100000101001110010111011110001110001001111100011000110101011101110010110111010010100111011000001101101001000100101000110001010101011010111000101010011010101011100001111000010100011010111110000101011100010100101101110110100011011010011001001000101101011111000110100010101100100001100000110111011110000000011100111000111110000001010001110001000110011000011011111100000010010010110010101011010110101010110110001011101001100110000000010111100010000111110101110001011000001001001111110110100000100101100101100010011010001111001001100101010100000110101101100010000000110100010011001100000000000101101100010101100101110101100001101000010010011011010001010010001010011110010100000111100100101111001000001101011001101010010000011011100111001010001010001000000111111010110000011110001001111011011110010101101000011100011110111110100010101101001111001101101001100011110001011001110011010101111011100101010111011001011101001000101100000001111011001010111001001101010000111001110111011110011011010111110000000001101101001100001101100100110001100011001100101001011011000100000010010011000010111111010001100111111000110100001000011010010100101010011001101000011011100000001001010101001111000000111001000101110000110001110111011011011100101100001000000000001000001111101011001100010111111011011100011010101011101010110101111110110000101000000010000111010000010000100111100000101100000001000101010110010101010110110000011010001110110110101010000101010010101000000101011010010111101111101011110001

`define PROTOTYPE_A_HIGH 2000'b00111011010010101000110100100010010110011110111001110100011000101111000111101010100111101010010010001111110001011111100001100100010101100111111100000100010100011101011100000000111011011011010101001010000100011100011110110000000101110100010010000111001101110011011100110000110001001101010011111011110100110101000001110111011100110001001101111000101100111111000001011001011111010011111010100000010001110010111010001000001101000110111011010111110001100110010101011110101101001111101011101111100011100100001101111000111111101100000001101110010111011110001110010101100111111001000101011101110010110111000010100110011000001101101010100101011000110001010101011000111000101010011001001011100001111000010100011010111110000101101100000100101101110110100011011010011001001000101101011000000110100001001100100101001000110111000010101010011100111000111100000001010001110001000110011000011011111100010110001110110010101011010110101000101010001011101001100110000010010111100010000111110001010001011001100101001111001110100000100101100101100010011010001111001001100101010000000110101101100010000000110100001100001100000011100101101100010101100101110001100001101000011010011011010001010011001100111110010100000111100100101111001000001101011001101010010000011011101011001010001010001000000111111010110011011011001001111011101110010101101000011100011110111110010010101101001111001101101001100011101101011001110011010100001011100101010111011011011101001000101101110011111011001010111001001001010000111001111011010000011011010111110000000001101101001100001010100100110001100011001100101001011011000100000010100011000010111111010001100111111000110100101000011010010100101010011001101000011101110000001001010101001111000000111001000001010001000000110111011011011100101100001000000000001000001111101011001100010111111011011100011010101011101010110101110110110000101000000010000111010000010100100111100000101100000001010110110110010101010110110000011010001110110110001010000101010010100110000101011010010111101111101011110000

`define PROTOTYPE_A_LOW 2000'b00111011010001110000110100100010010100011110111001110100011000101111000111101010100111101010010010001111110001011111100001100100010101100111111100110100010101101101011100000000000011011011010101001010000100001100011110110000000101110100010010000111001101110011011100110000101101001101010011111011110100110101000001110111011100110001100101111000101100111111001111011001010111010011111010100000010110110010111010001000001111000000111011010111110001100110010101011110101101001111101011101111100011100100001101111000111111101100000011101110010111011110001110001001111100111001000101011101110010110111000010100001011001001101101010100101001000110001011110101010111111101010011010101011100001111000010100011010111110000101001100010100010101110110100011011010011001001000100011011111000110111001001100100001110000110111011110011010011100111000111110000001010001110001000110011000011011111100000010000110110010101011010110100110110110001011101001100110000010010111100010000111110101110001011000010101001111000110100000100101100101100010011010001111001001100101010000000110101101100010000000110100010011101100000000000101101100010101100101101101100001101000010010011011010001010010001010000110010100000111100100101111001000001011011001101010010000011011110111001101001010001000000111111010110100011011111001111011101110010101101000011100011110111111010010101011001111001101101001100011101101011001110011010101111011100101010111011001011101001000101101101101111011001010111001010110010000111001111011011110011011010111110000000001101101001100001010100100110001100011001100101001011011000100000011010011000010111111010001100111111000110100010100011010010100101010011001101000011010110000001001010101001111100000111001000101110000110001110111011011011100101100001000000001001000001100001011001100010111111011011100011010101011101010110101111110110000101000000000000111010000010000100111100000101100000000100101010110010101010110110000011101001110110110001010000101010010101110000101011010010111101111101000001001

`endif

