`include "const.vh"

module associative_memory #(
	parameter AM_NUM_FOLDS, 
	parameter AM_NUM_FOLDS_WIDTH, 
	parameter AM_FOLD_WIDTH  
) (
	input						clk,
	input						rst,

	input						hvin_valid,
	output						hvin_ready,
	input	[`HV_DIMENSION-1:0]	hvin,

	output						dout_valid, 
	input						dout_ready,
	output reg					valence,
	output reg					arousal
);

	reg		[AM_FOLD_WIDTH-1:0]			similarity_hv;
	reg 	[`DISTANCE_WIDTH-1:0]		distance_p; 
	reg 	[`DISTANCE_WIDTH-1:0]		distance_n;   
	wire 	[`DISTANCE_WIDTH-1:0]		distance;

	wire 	hvin_fire;
	wire  	dout_fire;

	reg 	[AM_NUM_FOLDS_WIDTH-1:0] 	fold_counter;
	reg 	[2:0]						prototype_counter;

	// These need to be declared here to use the indexing method done for assigning to similarity_hv
	localparam PROTOTYPE_V_PLUS =   2000'b00111011010010110000110101010010010100111110111001110100011000101111000111101010100111101010010010001111110001011110100001100100010100010111111100100011001111001101011100011000111011011011010110010010000100100011111000110101100010001100101000110100011101111001000000000111101101011111010001100111111010110100101101110111100100110001000011111000101101001111001111011001010111010011111010100000010110001010111010100100000010000101100100001111101101110110011001011110101101000001100000100100101100101001001001001000110100110101110000101001100011000100001001001110111000100101100001010011110010110111010010100001011011101101101010100101000100110001011101101100111111101000001010101011100001111001100100111001111110111101101001111111110110011101100111000111100111010011110100001101010110011000110101011001100001110101010010100010011100111010101110000001010001110001000110011000011011111100000010001110110010101011010101001000110110110011101000000101110010010111100110101010010011111000001100111000100110111110111100010011100110111100101010001100101001110111001110011011101101100010000111110100010001110000000011100101101100010101100101001101100001101000010010001011010001010101000011100110010111111011100110110001101100101100110010110110001010000001010100100011001101101101100110011101011000100010111110111001110110010100100011111100011101010000011010101101001111001101101001100011101101011001110011010101111011100101001011010111000010101001100011001100111011110011001011110010100010111111101010011110101011010011101010100000100100110010011001100010001111100001011100011001100011111010000011010011011110111111010001100111111000110100001000011010000100101010011001101000011010110011010000100101001111000011100011010110110000000111000010010001001110001000011100111100110100010011110100011100101000101001011100000110100101101010110110011110110000101000000000000111010000010100100111100000101100000000110101010110010101010110110000011011111110110110110010000101010010100110000101011010010111101111101000000000;
	localparam PROTOTYPE_V_MIN  =   2000'b00111011010001110000110100100010010100011110111000010100011000101111000111101010100111101010010010001111110001011111100001100100010101100111111100000011001110101101011100011000000011011011010110010001100100100011111000110101100010001100100000111000011101111001000000000111101101011111010001101011011010110100101101110111100100110001110111111000101101001111001111011001010001010011111010100000010001110010111010110100010101000101100100001111101101110110011001011110101101001111010000100100101100101001011111001100110100110101110011001001110011000100001001001110111000000100010101010011110010110111001010100111011000001101101001000100101000110001011101011100111000101000001010001011100001111001100100000001111110111100001001111111010010011100000111000111111011010011010100001101010110001000110101011001000001110101001110100000011100111010101110000001010001110001000110011000011011111100000010010010110010101011010110101000110110110011101000000101110010010111100001101010011001111000001100111000100110111000111000010101111110111100101010001101001001101111010111100011101101100001100000110100010011110000000000000101101100010101100101110101100001101000010010011011010001010101000011100110010111111011100110110001101011101100110010110110001010000001010100100011001101101101100110011101010000100010111110111000000110010100100011111100011101010000011010101101001111001101101001100011110001011001110011010101111011100101000111010111000000101001100011011101111011110011001011110010100101111111101010011110101011010011101011010000100100110010011001100010001111100001011100101001000001000100000011010011011110111111010001100111111000110100001000011010010100101010011001101000011011100011101000100101001111000011111111010110110000110111000010010001001111001000011100111100110100010010100100111100101000101001011100000110100101101010110110011110110000101000000010000111010000010000100111100000101100000001000101010110010101010110110000011010001110110110101010000101010010101000000101011010010111101111101011110001;
	localparam PROTOTYPE_A_HIGH =   2000'b00111011010010101000110100100010010110011110111001110100011000101111000111101010100111101010010010001111110001011111100001100100010101100111111100000011001111011101011100011100111011011011010110010001100100100011111000110101100010001100101100111000011101111001000000000111101101011111010001101011111010110100101101110111100100110001001111111000101101001111000001011001011111010011111010100000010001110010111011100100010011000101100100101110101101110110011001011110101001000001000011010100101100101001010111001000110100110101110011001001110011000100001001001110111000001101100101010011110010110111010010100110011000001101101010100101011000110001011101011100111000101000001001001011100001111001100100110001111110111101111001111111110110011100000111000111111011010011000100001101010110000000110101011001000001110101001110100010011100111010101100000001010001110001000110011000011011111100010110001110110010101011010110101000110110110011101000000101110010010111100001101010011101111000001100111000100110111000110000010011011110111100101010001100101001110111110111011111101101100001100000110100010011110000000011100101101100010101100101110001100001101000011010011011010101010100000011100110010111111011100110110001101011101100110010110110001010000001010100100011001101101101100110011101010000100011111110111010000110010100100011111100011101010000011010101101001111001101101001100011101101011001110011010101111011100101010111010111000010101001100011011101111011110011001011110110100010111111101010011110101011010011101011000000100100110010011001100010001111100001011100101001011011111011000011010011011110111111010001100111111000110100101000011010010100101010011001101000011101110011010000100101001111000011100011010110110001000111000010010001001110111000011100111100110100010011100110111100101000101001011100000110100101101010110110011110110000101000000010000111010000010100100111100000101100000001010110110110010101010110110000011010001110110110001010000101010010100110000101011010010111101111101011110000;
	localparam PROTOTYPE_A_LOW  =   2000'b00111011010001110000110100100010010100011110111001110100011000101111000111101010100111101010010010001111110001011111100001100100010101100111111100110011001110101101011100011011000011011011001010010010000100100011111000110101100010001100101000100100011101111001000000000111101101011111010001101001011010110100101101110111100100110001101011111000100101001111001111011001010111010011111010100000010110001010111010110100010011000101100111001111101101110110011001011110101001001111100000100100101100101001011111001100110100110101110000101001110011000100001001001110111000100101100101010011110010110111010010100001011001001101101010100101001000110001011100101100111111101000001010101011100001111001100100110001111110111101111001111111010110011101100111000111100111010011110100001101010110011000110101011001101001110101010010100010011100111010101110000001010001110001000110011000011011111100000010000110110010101011010110101000110110110011101000000101110010010111100001101010010011111000001100111000100110110000111100010101100110111100101010001100101001110111101111101011101101100010000000110100010000010000000000000101101100010101100101101101100001101000010010011011010001010101001011100110010111111011100110110001101011101100110010110110001010000001010100100011001101101101100110011101010000100010111110111001110110010100100011111100011101010000011010101011001111001101101001100011101101011001110011010101111011100101001011010111000010101001100011011100111011110101001011110010100010111111101010011110101011010011101011110000110100110010011001100010001111100001011100101001100011000100000011010011011110111111010001100111111000110100010100011010010100101010011001101000011010110011101000100101001100000011101111010110110000110111000010010001001111001000011100111100110100010110101000111100101000101001011100000110100101101010110110011110110000101000000010000111010000010000100111100000101100000000100101010110010101010110110000011101001110110110001010000101010010101110000101011010010111101111101000001001;

	hv_binary_adder #(
		.AM_NUM_FOLDS          (AM_NUM_FOLDS),
		.AM_NUM_FOLDS_WIDTH    (AM_NUM_FOLDS_WIDTH),
		.AM_FOLD_WIDTH         (AM_FOLD_WIDTH)
    ) BIN_ADDER (
		.hv			(similarity_hv),
		.distance	(distance)
	);

	assign hvin_fire 	= hvin_valid && hvin_ready;
	assign hvin_ready	= prototype_counter == 0 && fold_counter == 0;

	assign dout_fire 	= dout_valid && dout_ready;
	assign dout_valid	= prototype_counter == 4;

	always @(posedge clk) begin
		if (rst || dout_fire)
			prototype_counter <= 0;
		else if (fold_counter == AM_NUM_FOLDS-1)
			prototype_counter <= prototype_counter + 1;
	end

	always @(posedge clk) begin
		if (rst || fold_counter == AM_NUM_FOLDS-1 || dout_fire)
			fold_counter <= 0;
		else if (hvin_fire || (fold_counter > 0 && fold_counter < AM_NUM_FOLDS-1) ||
				(fold_counter == 0 && prototype_counter > 0 && prototype_counter < 4))
			fold_counter <= fold_counter + 1;
	end

	always @(*) begin
		if (prototype_counter == 0) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_V_PLUS[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
		else if (prototype_counter == 1) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_V_MIN[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
		else if (prototype_counter == 2) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_A_HIGH[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
		else if (prototype_counter == 3) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_A_LOW[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
	end

	always @(posedge clk) begin
		if (prototype_counter == 0 || prototype_counter == 2) begin
			if (fold_counter == 0) 
				distance_p <= distance;
			else
				distance_p <= distance_p + distance;
		end		
	end

	always @(posedge clk) begin
		if (prototype_counter == 1 || prototype_counter == 3) begin
			if (fold_counter == 0) 
				distance_n <= distance;
			else
				distance_n <= distance_n + distance;
		end		
	end

	always @(posedge clk) begin
		if (prototype_counter == 1 && fold_counter == AM_NUM_FOLDS-1) begin
			valence <= distance_p >= (distance_n + distance);
		end

		if (prototype_counter == 3 && fold_counter == AM_NUM_FOLDS-1) begin
			arousal <= distance_p >= (distance_n + distance);
		end
	end

endmodule : associative_memory