`include "const.vh"

module associative_memory #(
	parameter NUM_FOLDS, 
	parameter NUM_FOLDS_WIDTH, 
	parameter FOLD_WIDTH  
) (
	input						clk,
	input						rst,

	input						hvin_valid,
	output						hvin_ready,
	input	[FOLD_WIDTH-1:0]	hvin,

	output						dout_valid, 
	input						dout_ready,
	output reg					valence,
	output reg					arousal
);

	reg   	[FOLD_WIDTH-1:0]		similarity_hv; 
	reg  	[`DISTANCE_WIDTH-1:0]	distance_vp;
	reg  	[`DISTANCE_WIDTH-1:0]	distance_vn; 
	reg  	[`DISTANCE_WIDTH-1:0]	distance_ap;
	reg  	[`DISTANCE_WIDTH-1:0]	distance_an;
	wire  	[`DISTANCE_WIDTH-1:0]	distance;

	reg 	[NUM_FOLDS_WIDTH-1:0] 	fold_counter; 
	reg 	[2:0]					prototype_counter;
  
	wire 	hvin_fire; 
	wire  	dout_fire;

	localparam PROTOTYPE_V_PLUS =   2000'b00111011011111000010011010001111111101001100011110000011001000001000101111100011111001001000000000001110110111011100111011100011011000001011110101100011100010101001110111111010011101100101100010011101011110011110010010111001010010110010110011101001010000001101101111010010010100011001110000100000010001001001101011001111100000011110100100100110000010101101001011011001011001001011001100011000110011011100100000100110000110000001011010010000001110011100111000101011100010010110011011111000011111010010101000110001110000110011001000010111001111100011001000001011100111001110010010011100000111100011111011100011101101011110101011001110011101111010111000011111100001000010110000010001001010110111110000111010110111010010000010111001110010111011010101100010100000000001110001011110110001101001101001111010010111010111011010100010000101000111010001001100011001111101100000100110010000011110011010100101001010000010101001011001100011101001110110111111101001011110001001000101000000011011110011000000100100010101100110010010101111110010111000111110001111000100010010011011010110001011000011011010000000011100111111001101101001110101010110111001111111101000101010001011101111101101100001101001010110010011100100101101101011001010100101110011010110100000011100101111110000010000100000000001110111101000100001101001010100111010010011010001101110100000010010110011100110101110001000100000100010110111011011100101110100101111110111000110101000100010000110110100011100001000001110100001110110010111010001111001001011010100001000101001011100101010001000110001111000101001001111001111111011101010111010110111100110110000100011011011001110011111010111110101000110101011100110000001001010001111110011111111010100001111010111000010001000011101001001011010101011001110111011101110011000001100001111110110101000111010000100011000100111011000011011000110010000000000100010011000011010100001100111111101110010000010010011101111110000110110011110100000001000110000110110000010001011011000101011110110010100000111001111001011;
	localparam PROTOTYPE_V_MIN  =   2000'b00111010011111000010011011111111111101111100011110000011001000001000101111100011111001001000000010100110110111011100111010100011010000001011110101110011100010101001110111111010011101100101100010011101011110011110000110111001000010100010001111101001010000001100101111010110010100001001110000100111100001001001101010111111100010011110100100100110000010101101001011011001011001001011001100011000110011011100100000100110000110010011011010010000010001011100111000101011100010010110011001111000011111010001111000100001110000110011001000010011001111100011001000101000000111001111100110011100000111010011111011100011101101011111101010111110011001111010111000011111100001000010110000010001000000010111110000111010110111010010000010111001110011001011010101111010001100000001110001011110110001000010101001110101010100110111011010101100000101000111011011001100011001111110000000100110010000011110000110100101001010111010101001011001100011101001110110111111010000101110001001000001000000011011110011011000100100010011100110010010101111110010111001111110001111000101011110011011010110001011000011011010000000011100111111001101101001110101010110111001111111101000101010001011101111101101100001101001010001010011100100101010101011001010100101110000010110100000011100101111110000001111000000000011010111101000100001101010100000011000010011010001101110100100010010110011100110001110001000100000100010110110111100100101110100100111110110110111011000100010000110110100011010100000000000100001110110010111011001111001011010110100001000101000000010101010001010010001111001011001001111001111111011110110111010110111100110110011000011011011001110011110010111110111100110110011100110001101001010001001110011111111010100001100010111000010001000011101001001011010101011001110111000001110011000001100001111110110101000111010000100011000100101100000011011000110100000110000100100100100011010100001100111111101110010000010010011101111110000110110011001111000000110110011110110000010001011011000101011110110010100000111001111001011;
	localparam PROTOTYPE_A_HIGH =   2000'b00111001111111000010011010111111111100001100011110000011001000001000101111100011111001001000000010000110110110011100111010100011011000001011110101101111100010101001110111111010011101100101100010011101011110011110011010111001001010110010110011101001010000001101101111010110010100001001110000100011100001001001101010001111100001011110100100100110000010101101001011011001011001001011001100011000110011011100100000100110000110001111011010010000001001011100111000101011100010010110011010011000011111010001010000100001110000110011001000010111001111100011001010001011100111001111100110011100000111111011111011100011101101011100101011001110011101111010111000011111100001000010110000010001000101110111110000111010110111010010000010111001110011001011010101100010011000000001110001011110110001010001111001111101010111110111011010100010000101000111011011001100011001111110000000100110010000011110011010100101001010111010101001011001100011101001110110111111101000011110001001000101000000011011110011111000100100010011100111010010101111110010111000111110001111000100011110011011010110001011000011011010000000011100111111001101101001110101010110111001111111101000101010001011101111101101100001101001010101010000000100101010101011001010100101110011010110100000111100101111110000000011000000000011110111101000100001101110010100011110010011010001101110100000010010110011100110101110001000100000100010110110101111100101110100100111110110110111101000100010000110110100011110001000001010100001110110010111011101111001011010110100001000101000011110101010001010011111111000101001001111001111111011101010111010110111100110110000100011011011001110011101110111001111100110110011100110011101001010000111110011111111010100001100010111000010001000011111001001011010101011001110111000001110011000001100001111110110101000111010000100011000100111011000011011011011010000110000100001000000011010100001100111111010110010000110010011101111110000110110011001111000000110110111110110000010001011011000101011110110010100000111001111001011;
	localparam PROTOTYPE_A_LOW  =   2000'b00111011011111000010011010001111111101001100011110000011001000001000101111100011111001001000000001001110110111011100111010100011011000001011110101110011100010101001110111111010011101100101100010011101011110011110001010111001010010110010001111101001010000001100101111010110010100011001110000001001100001001001101011111111100000011110100100100111110010101101011011011001011001001011001100011000110011011100100000100110000110000111100010010001111010011100111000101011100010010110011011111000011111010010111000110001110000110011001000010111001111100011001001101011100111001110010110011100000111011011111011100011101101011110101010111110011101111010111000011111100001000010110000010001001000110101110000111010110111010010000010111001110010111011010101100010100000000001110001011110110001100111101001110100010100110111011010100010000101000111011111001100011001111101100000100110010000011110001110111101001010000010101001011001100011011001110110111111010001111110001001000101000000011011110011000000100100011011100111010010101111110010111000111110001111000100101110011011010110001011000011011010000000011100111111001101101001110101010110111001111111101000101010001011101111101101100101101001001001010011100100101101101011001101100101110011010110100000011100101111110000001100100000000011110111101000100001101101010100011001010011010001100000100010010010110011100110001110001000100000100010110110111110100101110100101001110111000111011000100010000110110100011100111000000000100001110110010111011001111001001010110100001100101001111110101010001001110001111000101001001111001111111011101010111010110111100110110000100011011011001110011110010111110100010110110011100000000001001010001001110011111111010100001100010111000010001000011101001001011010101011001110111000001110011000001100001111110000101000111010000100011000100111011000011011000110000000110000100000111000011010100001100111111101110010000110010011101111110000110110011110111000000110110011110110000010001011011000101011110110010100000111001111001011;	

	assign hvin_fire 	= hvin_valid && hvin_ready;
	assign hvin_ready 	= prototype_counter == 0;

	assign dout_fire 	= dout_valid && dout_ready;
	assign dout_valid 	= prototype_counter == 4 && fold_counter == 0;

	always @(posedge clk) begin
		if (rst || dout_fire)
			fold_counter <= NUM_FOLDS-1;
		else if (prototype_counter == 4 && fold_counter != 0) 
			fold_counter <= fold_counter - 1;
	end

	always @(posedge clk) begin
		if (rst || (prototype_counter == 4 && fold_counter != 0) || dout_fire) 
			prototype_counter <= 0;
		else if (hvin_fire || (prototype_counter > 0 && prototype_counter < 4))
			prototype_counter <= prototype_counter + 1;
	end

	hv_binary_adder #(
		.NUM_FOLDS          (NUM_FOLDS),
		.NUM_FOLDS_WIDTH    (NUM_FOLDS_WIDTH),
		.FOLD_WIDTH         (FOLD_WIDTH)
    ) BIN_ADDER (
		.hv			(similarity_hv),
		.distance	(distance)
	);

	always @(*) begin
		if (prototype_counter == 0) begin
			similarity_hv = hvin ^ PROTOTYPE_V_PLUS[(fold_counter * FOLD_WIDTH) +: FOLD_WIDTH];
		end
		else if (prototype_counter == 1) begin
			similarity_hv = hvin ^ PROTOTYPE_V_MIN[(fold_counter * FOLD_WIDTH) +: FOLD_WIDTH];
		end
		else if (prototype_counter == 2) begin
			similarity_hv = hvin ^ PROTOTYPE_A_HIGH[(fold_counter * FOLD_WIDTH) +: FOLD_WIDTH];
		end
		else if (prototype_counter == 3) begin
			similarity_hv = hvin ^ PROTOTYPE_A_LOW[(fold_counter * FOLD_WIDTH) +: FOLD_WIDTH];
		end
	end

	always @(posedge clk) begin
		if (prototype_counter == 0 && hvin_valid) begin
			if (fold_counter == NUM_FOLDS-1)
				distance_vp <= distance;
			else
				distance_vp <= distance_vp + distance;
		end

		if (prototype_counter == 1) begin
			if (fold_counter == NUM_FOLDS-1)
				distance_vn <= distance;
			else
				distance_vn <= distance_vn + distance;
		end

		if (prototype_counter == 2) begin
			if (fold_counter == NUM_FOLDS-1)
				distance_ap <= distance;
			else
				distance_ap <= distance_ap + distance;
		end

		if (prototype_counter == 3) begin
			if (fold_counter == NUM_FOLDS-1)
				distance_an <= distance;
			else
				distance_an <= distance_an + distance;
		end
	end

	always @(posedge clk) begin
		if (fold_counter == 0 && prototype_counter == 1) 
			valence <= distance_vp >= (distance_vn + distance);

		if (fold_counter == 0 && prototype_counter == 3)
			arousal <= distance_ap >= (distance_an + distance);
	end

endmodule : associative_memory
