`include "const.vh"

module associative_memory #(
	parameter AM_NUM_FOLDS, 
	parameter AM_NUM_FOLDS_WIDTH, 
	parameter AM_FOLD_WIDTH  
) (
	input						clk,
	input						rst,

	input						hvin_valid,
	output						hvin_ready,
	input	[`HV_DIMENSION-1:0]	hvin,
 
	output						dout_valid,  
	input						dout_ready,
	output reg					valence,
	output reg					arousal
);

	reg		[AM_FOLD_WIDTH-1:0]			similarity_hv;
	reg 	[`DISTANCE_WIDTH-1:0]		distance_p; 
	reg 	[`DISTANCE_WIDTH-1:0]		distance_n;   
	wire 	[`DISTANCE_WIDTH-1:0]		distance;
   
	wire 	hvin_fire;
	wire  	dout_fire;

	reg 	[AM_NUM_FOLDS_WIDTH-1:0] 	fold_counter;
	reg 	[2:0]						prototype_counter;

	// These need to be declared here to use the indexing method done for assigning to similarity_hv
	localparam PROTOTYPE_V_PLUS =   2000'b00011011110010010000101010110001111100000011111000011101010000011111100000010111111110000101100011001111101111000010001100100100110111010111111111010100010110000001011110001111111010100101001010010011100001110110011001101010101010000101011010001110110101101110000101100111111000001011001101001000001100111010101001011110001111110100010110001100010010101010111000111010110100111110000101111000001010101001000010010110000111110101100100101111000111100110001010000001100001110101000101101000000011010111000100110110001110011100100101001111000101111010111111111110001001010001101101101011101101011000100111101000110100101100011001000110011100010110000011000001000110110111100111000101100000110011011010010101001000001100001111011111011000100010101100110110000001001001101110110001110010110000101100001001001001011100001111000000000010111001000001100001001101100100011010001000110001110001100000010000111100101010000110110111110101110000010001010001101110010100001100001001110110110000101100001101110001001110100010010011100010000000010111111000101101101000000001011110001110000001100101100011001000110100000001110011000000011001101010000010001110111111000110011000111110111000000100100101000000011111100000111111110000010011010100001011010001111011010000101011011000100100000000111101111000000011001110100100010101110101001100101100010000111011011010110110001000001001110010011000111110010000111101101100100110100101001011111011100010111101010110010011111110101111001101011111100100010101011001001110010000101111101110000010001001101000010101111111001101000010001011001011000111000000111111010100000011011111010000010000000011010111101000111110010101011100100101011101111101010100101001011100000000000011100100110101010101111101010110111110111100101010010000010011100000100110111010010100010000010001000011011100100011100100111010001110110100011010000001010000001101100011000110010000110000000001011100010001011001110101101011010100100001111100001101100010111101011110001010110111100000111010110000001100;
	localparam PROTOTYPE_V_MIN  =   2000'b00011011110010010000101010110001111101100011111011111101010000011111100000010111111110000001100011000111111111000010001100010100110111010111111111010100010111110001011110001110000010100101001010010011100001001001011001101010101010001101011011001110110000001011000101100101000100001011001101001000001111111010110111101110001111110111010110001100011110101010111100111010110010111110000100011000001010100101000010010110000000110101100100101111000100100110001010000001100001110100000101101000000011010111000100110110110110011100101011001111000001111010111000111110000101010001101101000011101101011000101111011100110100001100010100000110010000010110000011000001000110110111100101000101100110011111011010010101001000001100001111011111000100100010101110010110000001110101101110011001110010110000101100001001010110011100001111001110000010111001000011100001001101100100011010001000110001110001100000011100111100101010000001110111110101110000000001010001101110110110001100001100110100110000101101111101111001001110111011100011101110000000010000111001011101101000000001000110001110000000000010100011001000110000000001110000000000011001101010000010001110111111011110011000111010111000000100000111100000011111100110111111110100010011010010001011010001111011010000101011011000100100000000100110110000000011011010100000000110010101001100100100010000111000011010101010000000001001110010011110111111010000101101101100100110100101000111110001100010111101010111100111111110101111001101011110100000010101010001001111111001001111101010110010001001101000010101111111001101000010001011001011001011000000111111010100000011110111010000010000000011010111101000111110010101011100100000101101111101101100111101000100000000000000000101110111010101111101010111111110111100101010010100010011100000100110111010010100010000010000101011011100100011100100111010001110110100011010000000010000001101100011000110010111110000000111001100010000101001110101101011010100010001111100110101100011111101010000001010110111100000111010110100101100;
	localparam PROTOTYPE_A_HIGH =   2000'b00011011110010010000101010110001001111110011111000011101010000011111100000010111111110000001100011000111111111000010001100011100110111010111011111010100010111100001011110001111011010100101001010010011100001000001011001101010101010000101011011001110101001101110000101100111000100001011001101001000001011100110110101111110110111110111010110001100001110101010111100111010111100111110000101111000001010101001000000110110000000110101100100101111000111100110001010000001100001110101000101101000000011010111000100110110001110011100101111001111000010111010111011111110000110010001101101101011111101011000100110001100110100001100011001000110001100010110000011000001000110110111100101000101101011011111011010010101001000001101111111011111000100100001001100010110000001010101101110011001110010110000101100001001001001011100001111000000000010111001001101110101001101100100011010001000110001110001100000011100111100101010000001110111110101110000010001010001101110010111101100001001110110110000101101111101110111001110111001100011111110000000010000111001011101101000000001100110001110000010000101100011001000110000111001110011000000011001101010000010001110111111000110011000100010111000000100011111100000011111100000111111110100010011010100001011010001111011010000101011011000100100000000100101110000000011000010100110110111110101001100100100010000111000101010101010000100001001110010011111111110100000111101101100100110100101011011111101100010111101010110010111111110101111001101011110100100010101010001001110011001001111101101110010001001101000010101111111001101000010001011110011000111011100111111010100000011110111010000010000000011010111101000111110010101011100110101011101111101010100001101010100000000000011100001110101010101111101010110111110111100101010010000011011100000100110111010010100010000010001101011011100011011100100111010001110110100011010000001110000001101100011000100010111110000000001001100010000111001110101101011010100010001111100001101100011111001011110001010110111100000111010110000001100;
	localparam PROTOTYPE_A_LOW  =   2000'b00011011110010010000101010110001111101100011111011111010010000011111100000010111111110011101100010001111111111000010001100010100110111010111111111010100010110010001011110001111100010100101001010010011100001000110011001101010101010010101011001001110110101101110000101100011100101111011001101001010001100111010100011001110001111110111010110001100101110101010111010111010110010111110000111111000001010101101000010010110000111110101100100101111000111100110001010000001100001110101000101101000000011010111000100110110001110011100100111001111000101111010111111111110000111010001101101011011101101011000100111101100110101001100011101000110010000010110000011000001000110110111100100100101100000100011011010010101001000001100001111011111000100100010101100110110000001110101101110110011110010110000101100001001001100011100001111000000000010111001000011100001001101100100011010001000110001110001100000011010110100101010000110110111110101110000010001010001101110010100001100001001110110110000101101111101111001001110110011100011100010000000010111111000101101101000000001011110001110000001100101100011010100110000000001110011000000011001101010011110001110111111000110011000111110111000000100100100000000011111100110111111110101011011010010001011010001111011010000101011011000100100000000110110110000010011001110100111110100010101001100100100010000111111011010110110001000001001110010011000111111010000101101101100100110100101001011110011100010111101010110010111111110101111001101011110100000010101010001001111111000111111101001000010001001101000010101111111001101000010001011001011001111000000111111010100000011001111010000010000000011010111101000111110010101011100101101011101111101011100101001011100000000000011111101110101010101111101010110111110111100101010011100010011100000100110111010010100010000010001010011011100100011100100111010001110110100011010000000010000001101100011000110010000110000000001111100010001001001110101101011010000010001111100010101100010111111010010001010110111100000111010110001101100;
 
	hv_binary_adder #(
		.AM_NUM_FOLDS          (AM_NUM_FOLDS),
		.AM_NUM_FOLDS_WIDTH    (AM_NUM_FOLDS_WIDTH), 
		.AM_FOLD_WIDTH         (AM_FOLD_WIDTH) 
    ) BIN_ADDER (
		.hv			(similarity_hv),
		.distance	(distance)
	);

	assign hvin_fire 	= hvin_valid && hvin_ready;
	assign hvin_ready	= prototype_counter == 0 && fold_counter == 0;

	assign dout_fire 	= dout_valid && dout_ready;
	assign dout_valid	= prototype_counter == 4;
 
	always @(posedge clk) begin
		if (rst || dout_fire)
			prototype_counter <= 0;
		else if (fold_counter == AM_NUM_FOLDS-1)
			prototype_counter <= prototype_counter + 1;
	end

	always @(posedge clk) begin
		if (rst || fold_counter == AM_NUM_FOLDS-1 || dout_fire)
			fold_counter <= 0;
		else if (hvin_fire || (fold_counter > 0 && fold_counter < AM_NUM_FOLDS-1) ||
				(fold_counter == 0 && prototype_counter > 0 && prototype_counter < 4))
			fold_counter <= fold_counter + 1;
	end

	always @(*) begin
		if (prototype_counter == 0) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_V_PLUS[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
		else if (prototype_counter == 1) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_V_MIN[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
		else if (prototype_counter == 2) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_A_HIGH[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
		else if (prototype_counter == 3) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_A_LOW[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
	end

	always @(posedge clk) begin
		if (prototype_counter == 0 || prototype_counter == 2) begin
			if (fold_counter == 0) 
				distance_p <= distance;
			else
				distance_p <= distance_p + distance;
		end		
	end

	always @(posedge clk) begin
		if (prototype_counter == 1 || prototype_counter == 3) begin
			if (fold_counter == 0) 
				distance_n <= distance;
			else
				distance_n <= distance_n + distance;
		end		
	end

	always @(posedge clk) begin
		if (prototype_counter == 1 && fold_counter == AM_NUM_FOLDS-1) begin
			valence <= distance_p >= (distance_n + distance);
		end

		if (prototype_counter == 3 && fold_counter == AM_NUM_FOLDS-1) begin
			arousal <= distance_p >= (distance_n + distance);
		end
	end

endmodule : associative_memory