`include "const.vh"

module associative_memory #(
	parameter AM_NUM_FOLDS, 
	parameter AM_NUM_FOLDS_WIDTH, 
	parameter AM_FOLD_WIDTH  
) (
	input						clk,
	input						rst,

	input						hvin_valid,
	output						hvin_ready,
	input	[`HV_DIMENSION-1:0]	hvin,
 
	output						dout_valid,  
	input						dout_ready,
	output reg					valence,
	output reg					arousal
);

	reg		[AM_FOLD_WIDTH-1:0]			similarity_hv;
	reg 	[`DISTANCE_WIDTH-1:0]		distance_p; 
	reg 	[`DISTANCE_WIDTH-1:0]		distance_n;   
	wire 	[`DISTANCE_WIDTH-1:0]		distance;
   
	wire 	hvin_fire;
	wire  	dout_fire;

	reg 	[AM_NUM_FOLDS_WIDTH-1:0] 	fold_counter;
	reg 	[2:0]						prototype_counter;

	// These need to be declared here as localparams to use the indexing method done for assigning to similarity_hv
	// // NUM_FOLDS 1
	// localparam PROTOTYPE_V_PLUS =   2000'b00010011001110100010101101010000110100101010011001110100000101100111010101110111000001110010011100110111000111000010010010111111101000001111011111010011010010001000000000010011010010100110101010010011111101001100000001000110101111100100110011100000100011001100100100110111010000000101010011111001010111011011000111001111111000110001101000010011101111001100101100111001011000011000011110000000001010000100100111111101010100000101101101101010000001111001110111001110101110100001110111010110100000110011010001101010110001010100000101010011110110011000110001010010100100111101111010010111101110111010100010100000110100111100011001100110001110001001100011000110010100110100001011011011111100001000000110011101111110111011100011100011100011001001011100011001010011111101111011011110001000011011010010001011001110010000111101000011101100001010011010000001010010001110111010000110101100011101111100010010010110011101101101001111101010001011101000001011100000001100100010110010000010101110011000000111001110001101101010100011101110001100011011110010110101100000010010011101101010011100000100100110011011010000000011011110010000011001101001000011001111000010001111101011010000011011001001000000110010100011100110101110101000110111000110010001010001000101111110011110001011100000001111110000011011111011101000011011011101101001101111100100011110111000011010111110000011100011010100010111111000000010111100111001100111111001000100001000111110010000011011110011101000111000110101110000010000011101111111100000011111101011001100101101100001001100010110011101100011100101110011111011011000100001010010011011100110000001100000010111100101011011101000111101001100101101001001100101110111000000100011110000000000101100111111111111001010101100010010100110010110010111110110010100111011010010100111001111010000111000111100011110110111100100000100000000110011111110011001010000001101100000100011111011010000111100011110010111011101010110111101100000111110111000001111011110111101111001001101010010001100111000001010000000;
	// localparam PROTOTYPE_V_MIN  =   2000'b01010011000010100010101101010000110100101010011001110100000101100111010101110111000001110010011100001111100111000010110010111111101000001100011111010011010010001010100000010011110010100110101010010000011101001101100001000110101111110100111001111100100011001100000100110000001011000101010011110000010111011011010011001111111000110001101000010010101111001100101100111001011000011000011100000000001010000100000111111101011010000101101010101011010001111001110111001110101110100001110111011000100000110011000111101010110001010100000101010011110110011000110001010101100111011101111101010100101110111010110010100000110101111100011000000110011110001001100100000110010100110100010111011011111100001000000110011101111110111010000011100010010011001010111100011001010011111101111011011000001000011010010010001011000000010000111101000011101100001010011001000001010010001110111010000110101100011101111000010010101110010001101110101111110110001011101000001011100000001100100010110010000110101110011000001000101110001101101010100011101110001100011100110000100101000000010010011101101010010100111100100110011011010100000011011110010000011001101001000011001111000010001111101011011100011011001001000000110001100011100110101110101111110111001000010001101000100100001110011110001011100011000001111000011011111111001000011111010000010100011111100100011110110010011010111110000011100011010100101111111000000010111100111001100111111001000101001001011110010000011010000011101000111000110101100000010000011101111111101010011100001011001100101101110011001100010001011101100011100101110011111011011110100001010010011011100110010001000000010111100101011000001000111101001100101101000001100101111011000110011011001000111001101100111111111111001010011100010010100101110111100111110110010100111011101010100111001100110001001000111100011010110111100100000100000000110011111110011011010111001101100000100011111011010000111100011110010111011101010110111100100000111110100100001111011101111101111001001101010010001100111000001010000010;
	// localparam PROTOTYPE_A_HIGH =   2000'b01110010110000100010101101010000110100110010011001110100000101100111010101110111000001110010011101011111001111000010010010111111101000001111011111010011010010001010100000010011110010100110101010010010011101001110000001000110101111100100110011100111100011001100000100110111001000000101010011010000110111011011001011010111111000110001101000010011101111001100101100111001011000011000000010000000001010000100100111111101011010000101101101101011010000111001110111001110101110100001110111011000100000110011110001101010110001010100000101010011110110011000110001010010100101011101111010110100101110111010110010100000110101111100011001000110001110001001100100000110010100110100001011011011111100001000010110011101111110111100100011100010010011001011011100011001010000011101111010011000001000011010110010001011000000010000111101000011101100001010011010000001010010001110111010000110101100011101100000010010011110010011101101001111101010001011101000001011100000001100100010101110000110101110011000001001001110001101101010100011101110001100011011110001010101100000010010100101101010011100111100100110011011010000000011011110010000011001101001011011001111000010001111101011011110011011001001000000110011100011100110101110101111110111000110010011010000110100001110011110001011100011001111111000011011111011001000011111010011110100011111100100011110111010011010111110000011100011010100010111111000000010111100111001100111111001000011001000111110010000011011110011101000111000110101111100010000011101111111100000011111001011001100101101111101001100010110011101100011100101110011111011010110100001010010011011100110000001100000010111100101011011101000111101001100101101000101100101111011000000101011001000111001101100111111111111001010101100010010100101110111100111110110010100111011101010100111001000110001001000111100011111110111100100000101000000110011111110011010110111001101100000100011111011010000111100011110010111011101010110111100100000111110100100001111011101111101111001001101010010001100111000001010000010;
	// localparam PROTOTYPE_A_LOW  =   2000'b10010011001110100010101101010000110100101010011001110100000101100111010101110111000001110010011100010111000111000010110010111111101000001100111111010011010010001001000000010011110010100110101010010011111101001101100001000110101111100100110011100000100011001100100100110111010011000101010011101001010111011011010111001111111000110001101000010011001111001100101100111001011000011000011100000111001010000100100111111101010100000101101101101011000001111001110111001110101111100001110111010110100000110011011001101010110001010100000101010011110110011000110001010010100111011101111010001011101110111010110000100000110101111100011001000110001110001001100011000110010100110100001011011011111100010000000110011101111110111010100011100011100011001010111100011001001011111101111011011111001000011011010010001011001000010000111101000011101100001010011001000001010010001110111010000110101100011101111100010010101110011101101101001111111110001011101000001011100000001100100010110010010110101110011000000111001110001101101010100011101110001100011011110001100101110000010010011101101010011010000100100110000111010010000011011110010000011001101001000011001111000010001111101011010000011011001001000000110001100011100110101110101111110111001000011101110000000100001110011110001011100100000011111000011011111011001000011111011100001001101111100100011110110000011010111110000011100011010100000111111000000010111100111001100111111001000100001001011110010000011011110011101000111000110101111100010000011101111111100000011111101011001100101101100001001100010110011101100011100101110011111011011000100001010010011011100110000001110000010111100101011000001000111101001100111101011101100101110001000110011011110000000010001100111110111111001010101100010010100110010110010111110110010100111011010010100111001011110000111000111100011010110111100100100100000000110011111110011011010000001101100000100011111011010000111100011110010111011101010110111101100000111110111000001111011110111101111001001101010010001100111000001010000010;
	// // NUM_FOLDS 2
	// localparam PROTOTYPE_V_PLUS =   2000'b01110110001100010011001111110011111111101110011010010100010110001101011010000100001000111000010011100011110010100000111001000101110110001111011111101011010001010010100000101111110010100110101010010011111101110100000001000110101111100100110011100000100011001100100100110111010000000101010011111001010111011011000111001111111000110001101000010011101111001100101100111001011000011000011110000000001010000100100111111101010100000101101101101010000001111001110111001110101110100001110111010110100000110011010001101010110001010100000101010011110110011000110001010010100100111101111010010111101110111010100010100000110100111100011001100110001110001001100011000110010100110100001011011011111100001000000110011101111110111011100011100011100011001001011100011001010011111101111011011110001000011011011101010001011010001100111101011111101101111010000100011001010101010010100110011100011100000000000010010010011111011101011100000101111001101100000000011001101101110111110000001011101001101000011011001011011100000111100110011011011110111111100110100101111101010011001111111110101110111100001100101101110101100101011011001110011011011010001001111010101110100010001110011000110000011100110001011100111110100000011010101110101000110111000110010001010001000101111110011110001011100000001111110000011011111011101000011011011101101001101111100100011110111000011010111110000011100011010100010111111000000010111100111001100111111001000100001000111110010000011011110011101000111000110101110000010000011101111111100000011111101011001100101101100001001100010110011101100011100101110011111011011000100001010010011011100110000001100000010111100101011011101000111101001100101101001001100101110111000000100011110000000000101100111111111111001010101100010010100110010110010111110110010100111011010010100111001111010010000100111100011010110111101010000101001110110011011010000000010001111110000000011110010000111110000011010010111101101010100101101101111100101101000011001011110101010001001000100001011001110000110000111011111001;
	// localparam PROTOTYPE_V_MIN  =   2000'b01110110001100010011001111110011111111101110011010010011011110001101011010000100001000111000010011100001110010100010011001000101110110001100011111101011110001010010100000110111110010100110101010010000011101010101100001000110101111110100111001111100100011001100000100110000001011000101010011110000010111011011010011001111111000110001101000010010101111001100101100111001011000011000011100000000001010000100000111111101011010000101101010101011010001111001110111001110101110100001110111011000100000110011000111101010110001010100000101010011110110011000110001010101100111011101111101010100101110111010110010100000110101111100011000000110011110001001100100000110010100110100010111011011111100001000000110011101111110111010000011100010010011001010111100011001010011111101111011011000001000011010011101010001000100001100111101011111101101111010000010011001010011001010100110011100011100000000000010010010101111011101011100000110000101101001001100011001101101110111110000001000101001101000011011101011011100000111100110000111011110111100000110100101111010010011001110001110101110110010001011010101110101100101011011001110011011011010001001111000001110100010001110011000111100011100110001011100111001100000011010101110101111110111001000010001101000100100001110011110001011100011000001111000011011111111001000011111010000010100011111100100011110110010011010111110000011100011010100101111111000000010111100111001100111111001000101001001011110010000011010000011101000111000110101100000010000011101111111101010011100001011001100101101110011001100010001011101100011100101110011111011011110100001010010011011100110010001000000010111100101011000001000111101001100101101000001100101111011000110011011001000111001101100111111111111001010011100010010100101110111100111110110010100111011101010100111001100110010110100111100011010110111101010000100001100110010101010000000010110111110000000010110000000111110000100010001011101101010101010101101111100101101000110001011110101001101001000100001011001110000010000111011110001;
	// localparam PROTOTYPE_A_HIGH =   2000'b01110110001100010011001111100011111110101110011010010011010010001101011010000100001000111000010011100011110010100011111001000101110110001111011111101011010001010010101100101011110010100110101010010010011101110110000001000110101111100100110011100111100011001100000100110111001000000101010011010000110111011011001011010111111000110001101000010011101111001100101100111001011000011000000010000000001010000100100111111101011010000101101101101011010000111001110111001110101110100001110111011000100000110011110001101010110001010100000101010011110110011000110001010010100101011101111010110100101110111010110010100000110101111100011001000110001110001001100100000110010100110100001011011011111100001000010110011101111110111100100011100010010011001011011100011001010000011101111010011000001000011010111101010001010100001100111101011111101101111010000100011001010101001111100110011100011100000000000010001110101111011101011100000111111001101011001100011110101101110111110000001011101111110100011011110011011100000110110110000111011110111100000110100101111010010011001111111110101110111100001100111101110101100101011011001110011011011010001001111001001110100010001110011000111100011100110001011100111111100000011010101110101111110111000110010011010000110100001110011110001011100011001111111000011011111011001000011111010011110100011111100100011110111010011010111110000011100011010100010111111000000010111100111001100111111001000011001000111110010000011011110011101000111000110101111100010000011101111111100000011111001011001100101101111101001100010110011101100011100101110011111011010110100001010010011011100110000001100000010111100101011011101000111101001100101101000101100101111011000000101011001000111001101100111111111111001010101100010010100101110111100111110110010100111011101010100111001000110010110100111100011011110111101010000101010010110011011010000000110110111110000000010100001100111110000011010001011101101010101100101101111100101101000011101011110101011101001000100001011001110001000000111011111001;
	// localparam PROTOTYPE_A_LOW  =   2000'b01110110001100010011001111110011111111101110011010010100011000001110111010000100001000111000010011100101110010100000111001000101110110001100111111101011010001010010100000101111110010100110101010010011111101110101100001000110101111100100110011100000100011001100100100110111010011000101010011101001010111011011010111001111111000110001101000010011001111001100101100111001011000011000011100000111001010000100100111111101010100000101101101101011000001111001110111001110101111100001110111010110100000110011011001101010110001010100000101010011110110011000110001010010100111011101111010001011101110111010110000100000110101111100011001000110001110001001100011000110010100110100001011011011111100010000000110011101111110111010100011100011100011001010111100011001001011111101111011011111001000011011011101101001010100001100111101011111101101111010000111011001011011010010100110011100011100000000000010010010101111011101011100000101100101101100001100011001101101110111110000001000101101101000011011111101011100000111100110000111011110111111000110100101111010010011001110011110101110111000001100101101110101100101011011001110011011011010001001111010101110100010001110011000110000011100110001011100111101100000011010101110101111110111001000011101110000000100001110011110001011100100000011111000011011111011001000011111011100001001101111100100011110110000011010111110000011100011010100000111111000000010111100111001100111111001000100001001011110010000011011110011101000111000110101111100010000011101111111100000011111101011001100101101100001001100010110011101100011100101110011111011011000100001010010011011100110000001110000010111100101011000001000111101001100111101011101100101110001000110011011110000000010001100111110111111001010101100010010100110010110010111110110010100111011010010100111001011110011000100111100011010110111101010100101001100110011011010000000010001111110000000011110010000111110000101010010111101101010100101101101111100101101010111001011110101011101001000100001011001110000110000111011111001;
	// // NUM_FOLDS 4
	// localparam PROTOTYPE_V_PLUS =   2000'b11001101001100011010100101001101110100000010011011101010101111011000110000101011101100110010001111000000110001011110010110011101001110010111011100110100010000011101100000101111001010100110101010101011111101110100000001000110101111100100110011100000100011001100100100110111010000000101010011110001010111011011000000110000111000101101101100110011100111100010110111011010110110011100111101100000110010110011110111011000111010000011010101100001111111111010010001000110001011010111000101000000001101000110111100111011011110110111111101111010111100011110011011100100001000011001100011100011101101100010110011001010000010101100100010111010100100000111100010111100100011110100001011010101100011101110110110100100001110000011100011100011100011001001011100011001010011111101111011011110001000011011010011110101011010010000111101011111101010000101011010000000100101000000011110011010001011100000000010011100110001001011101101110011011000110100000101110110010100111001010100110110000011000111110000100110101111110000100010001100101111111101111001000101000100011001001111110110100011011101000111110110000000011101100011000110110000100001101001101010101011111110001111101000110000100100001001100011001110100011100110101110101000110111000110010001010001000101111110011110001011100000001111110000011011111010010100100111011101110101101100000111110000110000100010100001011011100011010011101000010100101110110011100101100011111101010000001101111001000111011010101000000010010101101001111001110111100010000011001010101000111001011000010001110100011100101000100011100010101001011101101111011010111101000011110000111010000111010001100000000010101001101001001101110111000000011001100101100110001000100011110000000001100010111111111110101010101100010010100110010110010111110110010100111011010010100111001111010011011111111100011010110111101001000000100100101100011110000110010001111111110000011110010110110010111100010011001001000111000010010001101010001100000000011101111111001101011110011000111101011100000111110101010000;
	// localparam PROTOTYPE_V_MIN  =   2000'b11001101001100011010100101111101110100100010011011101010100001011000000000101011101100110010001111000000110001011110010110011101001110010001011100110100010001101101100000100111001010100110101010101000011101110101100001000110101111110100111001111100100011001100000100110000001011000101010011110000010111011011010110110000111000101101101100110010100101100010110001011010110000011100111101100000110011110011110111011000111010000011010010100001111111111000010001000110001011010111000111000000001101011010000100111011011110110111111010111010111100000010011011100111000100011001100011100010001101100010110011001010000100001100101100111010101000000111101011011100100011110100000111000101100011101110001110100100001110000010000011100010010011001010111100011001010011111101111011011000001000011010010011110101010100010000111101011111101010000101011001000000100011011101101110011010001011100000000010011100110001001011101101110111111000110100100100010110010100111001010100110110000011000111110001010110101110110001010000001100101111111101111001100101000100011001001111110110100011010011000000110110000000011101100011000001110000100001101001101010101011111110001111101111101100100100001001100010001001100011100110101110101111110111001000010001101000100100001110011110001011100011000001111000011011111110010100100111010000010101101100000111110000110000100010100001011011100011010011101000101101011100110011110001100011111101001001001101111001000110011010101001000010010101101001111001110110100010011011001010101001001001011011110001110100011101001111100011100010101000011100001111010010111101000011110000111010100111010001100000000010101010001001001101110111000100011001100101100110110000011011001000000001100010111111111111001010011100010010100101110111100111110110010100111011101010100111001100110010101111111100011010110111101001000000100100101100011110000111010001111111110000011110001010110010111100010011001000110110100011010001101010000010011100100101111111001001010000011000111101100100000111110110010000;
	// localparam PROTOTYPE_A_HIGH =   2000'b11001101001100011010100101001101110111100010011011101010101111011000000000101011101100110010001111000000110001011110010110011101001110010011011100110100010000011101100000101011001010100110101010101010011101110110000001000110101111100100110011100111100011001100000100110111001000000101010011010000110111011011001000110000111000101001101100110011100111100010110001011010111000011100101101100000110010110011110111011000111010000011010101100001111111111100010001000110001011010111000011000000001101000110111100111011011110110111111010111010111100011110011011100000001100011001100011100011101101100010110011001010000110001100100010111010110100000111100100111100100100110100001010100101101011101110001110100100001110000100100011100010010011001011011100011001010000011101111010011000001000011010110011110101010100010000111101011111101010000101011010000000100101011100101110011010001011100000000010011100110001001011101101110111011000110100100101110110010100111001010100110110000101000111110001010111001110110000100011001100101111111101111001000101000100011001001111110110100011011011000111110110000000011101100011000110110000100001101001110110101011111110001111101000101100100100101001100010001111100011100110101001101111110111000110010011010000110100001110011110001011100011001111111000011011111010010100100111010011110101101100000111110000110000100010100001011111100011010011101000101101011110110011110001100011111101000001001101111001000110111010101011000010010101101001111001110000100010011011001010101001001001011100010001110100011100101000100011100010101001011101101111000110111101000011110000111001100111010001100000000010101001000001001101110111000100011001100101100110000000101011001000000001100010111111111110101010101100010010100101110111100111110110010100111011101010100111001000110010101111111100011011110111101001011001100100101100011110000111010001111111110111011110110110110010111010010011001000110100000010010001101010001110011100011101111111001101011110011000111101100100011011110101010000;
	// localparam PROTOTYPE_A_LOW  =   2000'b11001101001100011010100100111101110100100010011011101010100001011001110000101011101100110010001111000000110001011110010110011101001110010100111100110100010000101101100000101111001010100110101010101011111101110101100001000110101111100100110011100000100011001100100100110111010011000101010011101001010111011011010000110000111000101101101100110011000111100010110011011010110110011100111101100110110100110011110111001000111010000011010101100001111111111011010001000110001011010111000100100000001101011010011100111011011110110111111010111010111010000010011011000000001100011001100011100010011101100010110001001010000011001100100110111010101000000111101011011100100011110100001011010101100001101110110110100100001110000010100011100011100011001010111100011001001011111101111011011111001000011011010011110101010000010000111101011111100110000101011001000000100011000000011110011010001011100000000010011100110001001011101101110011011000110111100101110110010100111001010100110110000011000111110000100110101111110000100010001100101111111101111010100101000100011001001111110110101111011011000111110110000000011101100011000110110000100001101001101010101011111110001111101000110000100100001001100010011101100011100110101110101111110111001000011101110000000100001110011110001011100100000011111000011011111010010100100111011100010101101100000111110000110000100010100001011011100011010011101000110100101110110011101101100011111101011000001101111001000111011010101011000010010101101001111001110111100010011011001010101010101001011100110001110100011101001000100011100010101001011101101111011110111101000011110000111010000111010001100000000010101010001001001101110111010100011001100101100110110000011011110000000001100010111110111101001010101100010010100110010110010111110110010100111011010010100111001011110011011111111100011010110111101001000000100100101100011110000111010001111111110000011110010010110010111100010011001001010111100011010001101010000100000000111101111111001010010000011000111101011100000111110000010000;
	// NUM_FOLDS 8	
	localparam PROTOTYPE_V_PLUS =   2000'b00011011110010010000101010110001111100000011111000011101010000011111100000010111111110000101100011001111101111000010001100100100110111010111111111010100010110000001011110001111111010100101001010010011100001110110011001101010101010000101011010001110110101101110000101100111111000001011001101001000001100111010101001011110001111110100010110001100010010101010111000111010110100111110000101111000001010101001000010010110000111110101100100101111000111100110001010000001100001110101000101101000000011010111000100110110001110011100100101001111000101111010111111111110001001010001101101101011101101011000100111101000110100101100011001000110011100010110000011000001000110110111100111000101100000110011011010010101001000001100001111011111011000100010101100110110000001001001101110110001110010110000101100001001001001011100001111000000000010111001000001100001001101100100011010001000110001110001100000010000111100101010000110110111110101110000010001010001101110010100001100001001110110110000101100001101110001001110100010010011100010000000010111111000101101101000000001011110001110000001100101100011001000110100000001110011000000011001101010000010001110111111000110011000111110111000000100100101000000011111100000111111110000010011010100001011010001111011010000101011011000100100000000111101111000000011001110100100010101110101001100101100010000111011011010110110001000001001110010011000111110010000111101101100100110100101001011111011100010111101010110010011111110101111001101011111100100010101011001001110010000101111101110000010001001101000010101111111001101000010001011001011000111000000111111010100000011011111010000010000000011010111101000111110010101011100100101011101111101010100101001011100000000000011100100110101010101111101010110111110111100101010010000010011100000100110111010010100010000010001000011011100100011100100111010001110110100011010000001010000001101100011000110010000110000000001011100010001011001110101101011010100100001111100001101100010111101011110001010110111100000111010110000001100;
	localparam PROTOTYPE_V_MIN  =   2000'b00011011110010010000101010110001111101100011111011111101010000011111100000010111111110000001100011000111111111000010001100010100110111010111111111010100010111110001011110001110000010100101001010010011100001001001011001101010101010001101011011001110110000001011000101100101000100001011001101001000001111111010110111101110001111110111010110001100011110101010111100111010110010111110000100011000001010100101000010010110000000110101100100101111000100100110001010000001100001110100000101101000000011010111000100110110110110011100101011001111000001111010111000111110000101010001101101000011101101011000101111011100110100001100010100000110010000010110000011000001000110110111100101000101100110011111011010010101001000001100001111011111000100100010101110010110000001110101101110011001110010110000101100001001010110011100001111001110000010111001000011100001001101100100011010001000110001110001100000011100111100101010000001110111110101110000000001010001101110110110001100001100110100110000101101111101111001001110111011100011101110000000010000111001011101101000000001000110001110000000000010100011001000110000000001110000000000011001101010000010001110111111011110011000111010111000000100000111100000011111100110111111110100010011010010001011010001111011010000101011011000100100000000100110110000000011011010100000000110010101001100100100010000111000011010101010000000001001110010011110111111010000101101101100100110100101000111110001100010111101010111100111111110101111001101011110100000010101010001001111111001001111101010110010001001101000010101111111001101000010001011001011001011000000111111010100000011110111010000010000000011010111101000111110010101011100100000101101111101101100111101000100000000000000000101110111010101111101010111111110111100101010010100010011100000100110111010010100010000010000101011011100100011100100111010001110110100011010000000010000001101100011000110010111110000000111001100010000101001110101101011010100010001111100110101100011111101010000001010110111100000111010110100101100;
	localparam PROTOTYPE_A_HIGH =   2000'b00011011110010010000101010110001001111110011111000011101010000011111100000010111111110000001100011000111111111000010001100011100110111010111011111010100010111100001011110001111011010100101001010010011100001000001011001101010101010000101011011001110101001101110000101100111000100001011001101001000001011100110110101111110110111110111010110001100001110101010111100111010111100111110000101111000001010101001000000110110000000110101100100101111000111100110001010000001100001110101000101101000000011010111000100110110001110011100101111001111000010111010111011111110000110010001101101101011111101011000100110001100110100001100011001000110001100010110000011000001000110110111100101000101101011011111011010010101001000001101111111011111000100100001001100010110000001010101101110011001110010110000101100001001001001011100001111000000000010111001001101110101001101100100011010001000110001110001100000011100111100101010000001110111110101110000010001010001101110010111101100001001110110110000101101111101110111001110111001100011111110000000010000111001011101101000000001100110001110000010000101100011001000110000111001110011000000011001101010000010001110111111000110011000100010111000000100011111100000011111100000111111110100010011010100001011010001111011010000101011011000100100000000100101110000000011000010100110110111110101001100100100010000111000101010101010000100001001110010011111111110100000111101101100100110100101011011111101100010111101010110010111111110101111001101011110100100010101010001001110011001001111101101110010001001101000010101111111001101000010001011110011000111011100111111010100000011110111010000010000000011010111101000111110010101011100110101011101111101010100001101010100000000000011100001110101010101111101010110111110111100101010010000011011100000100110111010010100010000010001101011011100011011100100111010001110110100011010000001110000001101100011000100010111110000000001001100010000111001110101101011010100010001111100001101100011111001011110001010110111100000111010110000001100;
	localparam PROTOTYPE_A_LOW  =   2000'b00011011110010010000101010110001111101100011111011111010010000011111100000010111111110011101100010001111111111000010001100010100110111010111111111010100010110010001011110001111100010100101001010010011100001000110011001101010101010010101011001001110110101101110000101100011100101111011001101001010001100111010100011001110001111110111010110001100101110101010111010111010110010111110000111111000001010101101000010010110000111110101100100101111000111100110001010000001100001110101000101101000000011010111000100110110001110011100100111001111000101111010111111111110000111010001101101011011101101011000100111101100110101001100011101000110010000010110000011000001000110110111100100100101100000100011011010010101001000001100001111011111000100100010101100110110000001110101101110110011110010110000101100001001001100011100001111000000000010111001000011100001001101100100011010001000110001110001100000011010110100101010000110110111110101110000010001010001101110010100001100001001110110110000101101111101111001001110110011100011100010000000010111111000101101101000000001011110001110000001100101100011010100110000000001110011000000011001101010011110001110111111000110011000111110111000000100100100000000011111100110111111110101011011010010001011010001111011010000101011011000100100000000110110110000010011001110100111110100010101001100100100010000111111011010110110001000001001110010011000111111010000101101101100100110100101001011110011100010111101010110010111111110101111001101011110100000010101010001001111111000111111101001000010001001101000010101111111001101000010001011001011001111000000111111010100000011001111010000010000000011010111101000111110010101011100101101011101111101011100101001011100000000000011111101110101010101111101010110111110111100101010011100010011100000100110111010010100010000010001010011011100100011100100111010001110110100011010000000010000001101100011000110010000110000000001111100010001001001110101101011010000010001111100010101100010111111010010001010110111100000111010110001101100;
 
	hv_binary_adder #(
		.AM_NUM_FOLDS          (AM_NUM_FOLDS),
		.AM_NUM_FOLDS_WIDTH    (AM_NUM_FOLDS_WIDTH), 
		.AM_FOLD_WIDTH         (AM_FOLD_WIDTH) 
    ) BIN_ADDER (
		.hv			(similarity_hv),
		.distance	(distance)
	);

	assign hvin_fire 	= hvin_valid && hvin_ready;
	assign hvin_ready	= prototype_counter == 0 && fold_counter == 0;

	assign dout_fire 	= dout_valid && dout_ready;
	assign dout_valid	= prototype_counter == 4;
 
	always @(posedge clk) begin
		if (rst || dout_fire)
			prototype_counter <= 0;
		else if (fold_counter == AM_NUM_FOLDS-1)
			prototype_counter <= prototype_counter + 1;
	end

	always @(posedge clk) begin
		if (rst || fold_counter == AM_NUM_FOLDS-1 || dout_fire)
			fold_counter <= 0;
		else if (hvin_fire || (fold_counter > 0 && fold_counter < AM_NUM_FOLDS-1) ||
				(fold_counter == 0 && prototype_counter > 0 && prototype_counter < 4))
			fold_counter <= fold_counter + 1;
	end

	always @(*) begin
		if (prototype_counter == 0) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_V_PLUS[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
		else if (prototype_counter == 1) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_V_MIN[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
		else if (prototype_counter == 2) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_A_HIGH[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
		else if (prototype_counter == 3) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_A_LOW[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
	end

	always @(posedge clk) begin
		if (prototype_counter == 0 || prototype_counter == 2) begin
			if (fold_counter == 0) 
				distance_p <= distance;
			else
				distance_p <= distance_p + distance;
		end		
	end

	always @(posedge clk) begin
		if (prototype_counter == 1 || prototype_counter == 3) begin
			if (fold_counter == 0) 
				distance_n <= distance;
			else
				distance_n <= distance_n + distance;
		end		
	end

	always @(posedge clk) begin
		if (prototype_counter == 1 && fold_counter == AM_NUM_FOLDS-1) begin
			valence <= distance_p >= (distance_n + distance);
		end

		if (prototype_counter == 3 && fold_counter == AM_NUM_FOLDS-1) begin
			arousal <= distance_p >= (distance_n + distance);
		end
	end

endmodule : associative_memory
