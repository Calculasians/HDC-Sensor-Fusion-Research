`include "const.vh"

module associative_memory #(
	parameter AM_NUM_FOLDS, 
	parameter AM_NUM_FOLDS_WIDTH, 
	parameter AM_FOLD_WIDTH  
) (
	input						clk,
	input						rst,

	input						hvin_valid,
	output						hvin_ready,
	input	[`HV_DIMENSION-1:0]	hvin,
 
	output						dout_valid,  
	input						dout_ready,
	output reg					valence,
	output reg					arousal
);

	reg		[AM_FOLD_WIDTH-1:0]			similarity_hv;
	reg 	[`DISTANCE_WIDTH-1:0]		distance_p; 
	reg 	[`DISTANCE_WIDTH-1:0]		distance_n;   
	wire 	[`DISTANCE_WIDTH-1:0]		distance;
   
	wire 	hvin_fire;
	wire  	dout_fire;

	reg 	[AM_NUM_FOLDS_WIDTH-1:0] 	fold_counter;
	reg 	[2:0]						prototype_counter;

	// These need to be declared here to use the indexing method done for assigning to similarity_hv
	localparam PROTOTYPE_V_PLUS =   2000'b11001101001100011010100101001101110100000010011011101010101111011000110000101011101100110010001111000000110001011110010110011101001110010111011100110100010000011101100000101111001010100110101010101011111101110100000001000110101111100100110011100000100011001100100100110111010000000101010011110001010111011011000000110000111000101101101100110011100111100010110111011010110110011100111101100000110010110011110111011000111010000011010101100001111111111010010001000110001011010111000101000000001101000110111100111011011110110111111101111010111100011110011011100100001000011001100011100011101101100010110011001010000010101100100010111010100100000111100010111100100011110100001011010101100011101110110110100100001110000011100011100011100011001001011100011001010011111101111011011110001000011011010011110101011010010000111101011111101010000101011010000000100101000000011110011010001011100000000010011100110001001011101101110011011000110100000101110110010100111001010100110110000011000111110000100110101111110000100010001100101111111101111001000101000100011001001111110110100011011101000111110110000000011101100011000110110000100001101001101010101011111110001111101000110000100100001001100011001110100011100110101110101000110111000110010001010001000101111110011110001011100000001111110000011011111010010100100111011101110101101100000111110000110000100010100001011011100011010011101000010100101110110011100101100011111101010000001101111001000111011010101000000010010101101001111001110111100010000011001010101000111001011000010001110100011100101000100011100010101001011101101111011010111101000011110000111010000111010001100000000010101001101001001101110111000000011001100101100110001000100011110000000001100010111111111110101010101100010010100110010110010111110110010100111011010010100111001111010011011111111100011010110111101001000000100100101100011110000110010001111111110000011110010110110010111100010011001001000111000010010001101010001100000000011101111111001101011110011000111101011100000111110101010000;
	localparam PROTOTYPE_V_MIN  =   2000'b11001101001100011010100101111101110100100010011011101010100001011000000000101011101100110010001111000000110001011110010110011101001110010001011100110100010001101101100000100111001010100110101010101000011101110101100001000110101111110100111001111100100011001100000100110000001011000101010011110000010111011011010110110000111000101101101100110010100101100010110001011010110000011100111101100000110011110011110111011000111010000011010010100001111111111000010001000110001011010111000111000000001101011010000100111011011110110111111010111010111100000010011011100111000100011001100011100010001101100010110011001010000100001100101100111010101000000111101011011100100011110100000111000101100011101110001110100100001110000010000011100010010011001010111100011001010011111101111011011000001000011010010011110101010100010000111101011111101010000101011001000000100011011101101110011010001011100000000010011100110001001011101101110111111000110100100100010110010100111001010100110110000011000111110001010110101110110001010000001100101111111101111001100101000100011001001111110110100011010011000000110110000000011101100011000001110000100001101001101010101011111110001111101111101100100100001001100010001001100011100110101110101111110111001000010001101000100100001110011110001011100011000001111000011011111110010100100111010000010101101100000111110000110000100010100001011011100011010011101000101101011100110011110001100011111101001001001101111001000110011010101001000010010101101001111001110110100010011011001010101001001001011011110001110100011101001111100011100010101000011100001111010010111101000011110000111010100111010001100000000010101010001001001101110111000100011001100101100110110000011011001000000001100010111111111111001010011100010010100101110111100111110110010100111011101010100111001100110010101111111100011010110111101001000000100100101100011110000111010001111111110000011110001010110010111100010011001000110110100011010001101010000010011100100101111111001001010000011000111101100100000111110110010000;
	localparam PROTOTYPE_A_HIGH =   2000'b11001101001100011010100101001101110111100010011011101010101111011000000000101011101100110010001111000000110001011110010110011101001110010011011100110100010000011101100000101011001010100110101010101010011101110110000001000110101111100100110011100111100011001100000100110111001000000101010011010000110111011011001000110000111000101001101100110011100111100010110001011010111000011100101101100000110010110011110111011000111010000011010101100001111111111100010001000110001011010111000011000000001101000110111100111011011110110111111010111010111100011110011011100000001100011001100011100011101101100010110011001010000110001100100010111010110100000111100100111100100100110100001010100101101011101110001110100100001110000100100011100010010011001011011100011001010000011101111010011000001000011010110011110101010100010000111101011111101010000101011010000000100101011100101110011010001011100000000010011100110001001011101101110111011000110100100101110110010100111001010100110110000101000111110001010111001110110000100011001100101111111101111001000101000100011001001111110110100011011011000111110110000000011101100011000110110000100001101001110110101011111110001111101000101100100100101001100010001111100011100110101001101111110111000110010011010000110100001110011110001011100011001111111000011011111010010100100111010011110101101100000111110000110000100010100001011111100011010011101000101101011110110011110001100011111101000001001101111001000110111010101011000010010101101001111001110000100010011011001010101001001001011100010001110100011100101000100011100010101001011101101111000110111101000011110000111001100111010001100000000010101001000001001101110111000100011001100101100110000000101011001000000001100010111111111110101010101100010010100101110111100111110110010100111011101010100111001000110010101111111100011011110111101001011001100100101100011110000111010001111111110111011110110110110010111010010011001000110100000010010001101010001110011100011101111111001101011110011000111101100100011011110101010000;
	localparam PROTOTYPE_A_LOW  =   2000'b11001101001100011010100100111101110100100010011011101010100001011001110000101011101100110010001111000000110001011110010110011101001110010100111100110100010000101101100000101111001010100110101010101011111101110101100001000110101111100100110011100000100011001100100100110111010011000101010011101001010111011011010000110000111000101101101100110011000111100010110011011010110110011100111101100110110100110011110111001000111010000011010101100001111111111011010001000110001011010111000100100000001101011010011100111011011110110111111010111010111010000010011011000000001100011001100011100010011101100010110001001010000011001100100110111010101000000111101011011100100011110100001011010101100001101110110110100100001110000010100011100011100011001010111100011001001011111101111011011111001000011011010011110101010000010000111101011111100110000101011001000000100011000000011110011010001011100000000010011100110001001011101101110011011000110111100101110110010100111001010100110110000011000111110000100110101111110000100010001100101111111101111010100101000100011001001111110110101111011011000111110110000000011101100011000110110000100001101001101010101011111110001111101000110000100100001001100010011101100011100110101110101111110111001000011101110000000100001110011110001011100100000011111000011011111010010100100111011100010101101100000111110000110000100010100001011011100011010011101000110100101110110011101101100011111101011000001101111001000111011010101011000010010101101001111001110111100010011011001010101010101001011100110001110100011101001000100011100010101001011101101111011110111101000011110000111010000111010001100000000010101010001001001101110111010100011001100101100110110000011011110000000001100010111110111101001010101100010010100110010110010111110110010100111011010010100111001011110011011111111100011010110111101001000000100100101100011110000111010001111111110000011110010010110010111100010011001001010111100011010001101010000100000000111101111111001010010000011000111101011100000111110000010000;
 
	hv_binary_adder #(
		.AM_NUM_FOLDS          (AM_NUM_FOLDS),
		.AM_NUM_FOLDS_WIDTH    (AM_NUM_FOLDS_WIDTH), 
		.AM_FOLD_WIDTH         (AM_FOLD_WIDTH) 
    ) BIN_ADDER (
		.hv			(similarity_hv),
		.distance	(distance)
	);

	assign hvin_fire 	= hvin_valid && hvin_ready;
	assign hvin_ready	= prototype_counter == 0 && fold_counter == 0;

	assign dout_fire 	= dout_valid && dout_ready;
	assign dout_valid	= prototype_counter == 4;
 
	always @(posedge clk) begin
		if (rst || dout_fire)
			prototype_counter <= 0;
		else if (fold_counter == AM_NUM_FOLDS-1)
			prototype_counter <= prototype_counter + 1;
	end

	always @(posedge clk) begin
		if (rst || fold_counter == AM_NUM_FOLDS-1 || dout_fire)
			fold_counter <= 0;
		else if (hvin_fire || (fold_counter > 0 && fold_counter < AM_NUM_FOLDS-1) ||
				(fold_counter == 0 && prototype_counter > 0 && prototype_counter < 4))
			fold_counter <= fold_counter + 1;
	end

	always @(*) begin
		if (prototype_counter == 0) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_V_PLUS[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
		else if (prototype_counter == 1) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_V_MIN[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
		else if (prototype_counter == 2) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_A_HIGH[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
		else if (prototype_counter == 3) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_A_LOW[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
	end

	always @(posedge clk) begin
		if (prototype_counter == 0 || prototype_counter == 2) begin
			if (fold_counter == 0) 
				distance_p <= distance;
			else
				distance_p <= distance_p + distance;
		end		
	end

	always @(posedge clk) begin
		if (prototype_counter == 1 || prototype_counter == 3) begin
			if (fold_counter == 0) 
				distance_n <= distance;
			else
				distance_n <= distance_n + distance;
		end		
	end

	always @(posedge clk) begin
		if (prototype_counter == 1 && fold_counter == AM_NUM_FOLDS-1) begin
			valence <= distance_p >= (distance_n + distance);
		end

		if (prototype_counter == 3 && fold_counter == AM_NUM_FOLDS-1) begin
			arousal <= distance_p >= (distance_n + distance);
		end
	end

endmodule : associative_memory
