`include "const.vh"

module associative_memory #(
	parameter AM_NUM_FOLDS, 
	parameter AM_NUM_FOLDS_WIDTH, 
	parameter AM_FOLD_WIDTH  
) (
	input						clk,
	input						rst,

	input						hvin_valid,
	output						hvin_ready,
	input	[`HV_DIMENSION-1:0]	hvin,
 
	output						dout_valid,  
	input						dout_ready,
	output reg					valence,
	output reg					arousal
);

	reg		[AM_FOLD_WIDTH-1:0]			similarity_hv;
	reg 	[`DISTANCE_WIDTH-1:0]		distance_p; 
	reg 	[`DISTANCE_WIDTH-1:0]		distance_n;   
	wire 	[`DISTANCE_WIDTH-1:0]		distance;
   
	wire 	hvin_fire;
	wire  	dout_fire;

	reg 	[AM_NUM_FOLDS_WIDTH-1:0] 	fold_counter;
	reg 	[2:0]						prototype_counter;

	// These need to be declared here to use the indexing method done for assigning to similarity_hv
	localparam PROTOTYPE_V_PLUS =   2000'b00010011001110100010101101010000110100101010011001110100000101100111010101110111000001110010011100110111000111000010010010111111101000001111011111010011010010001000000000010011010010100110101010010011111101001100000001000110101111100100110011100000100011001100100100110111010000000101010011111001010111011011000111001111111000110001101000010011101111001100101100111001011000011000011110000000001010000100100111111101010100000101101101101010000001111001110111001110101110100001110111010110100000110011010001101010110001010100000101010011110110011000110001010010100100111101111010010111101110111010100010100000110100111100011001100110001110001001100011000110010100110100001011011011111100001000000110011101111110111011100011100011100011001001011100011001010011111101111011011110001000011011010010001011001110010000111101000011101100001010011010000001010010001110111010000110101100011101111100010010010110011101101101001111101010001011101000001011100000001100100010110010000010101110011000000111001110001101101010100011101110001100011011110010110101100000010010011101101010011100000100100110011011010000000011011110010000011001101001000011001111000010001111101011010000011011001001000000110010100011100110101110101000110111000110010001010001000101111110011110001011100000001111110000011011111011101000011011011101101001101111100100011110111000011010111110000011100011010100010111111000000010111100111001100111111001000100001000111110010000011011110011101000111000110101110000010000011101111111100000011111101011001100101101100001001100010110011101100011100101110011111011011000100001010010011011100110000001100000010111100101011011101000111101001100101101001001100101110111000000100011110000000000101100111111111111001010101100010010100110010110010111110110010100111011010010100111001111010000111000111100011110110111100100000100000000110011111110011001010000001101100000100011111011010000111100011110010111011101010110111101100000111110111000001111011110111101111001001101010010001100111000001010000000;
	localparam PROTOTYPE_V_MIN  =   2000'b01010011000010100010101101010000110100101010011001110100000101100111010101110111000001110010011100001111100111000010110010111111101000001100011111010011010010001010100000010011110010100110101010010000011101001101100001000110101111110100111001111100100011001100000100110000001011000101010011110000010111011011010011001111111000110001101000010010101111001100101100111001011000011000011100000000001010000100000111111101011010000101101010101011010001111001110111001110101110100001110111011000100000110011000111101010110001010100000101010011110110011000110001010101100111011101111101010100101110111010110010100000110101111100011000000110011110001001100100000110010100110100010111011011111100001000000110011101111110111010000011100010010011001010111100011001010011111101111011011000001000011010010010001011000000010000111101000011101100001010011001000001010010001110111010000110101100011101111000010010101110010001101110101111110110001011101000001011100000001100100010110010000110101110011000001000101110001101101010100011101110001100011100110000100101000000010010011101101010010100111100100110011011010100000011011110010000011001101001000011001111000010001111101011011100011011001001000000110001100011100110101110101111110111001000010001101000100100001110011110001011100011000001111000011011111111001000011111010000010100011111100100011110110010011010111110000011100011010100101111111000000010111100111001100111111001000101001001011110010000011010000011101000111000110101100000010000011101111111101010011100001011001100101101110011001100010001011101100011100101110011111011011110100001010010011011100110010001000000010111100101011000001000111101001100101101000001100101111011000110011011001000111001101100111111111111001010011100010010100101110111100111110110010100111011101010100111001100110001001000111100011010110111100100000100000000110011111110011011010111001101100000100011111011010000111100011110010111011101010110111100100000111110100100001111011101111101111001001101010010001100111000001010000010;
	localparam PROTOTYPE_A_HIGH =   2000'b01110010110000100010101101010000110100110010011001110100000101100111010101110111000001110010011101011111001111000010010010111111101000001111011111010011010010001010100000010011110010100110101010010010011101001110000001000110101111100100110011100111100011001100000100110111001000000101010011010000110111011011001011010111111000110001101000010011101111001100101100111001011000011000000010000000001010000100100111111101011010000101101101101011010000111001110111001110101110100001110111011000100000110011110001101010110001010100000101010011110110011000110001010010100101011101111010110100101110111010110010100000110101111100011001000110001110001001100100000110010100110100001011011011111100001000010110011101111110111100100011100010010011001011011100011001010000011101111010011000001000011010110010001011000000010000111101000011101100001010011010000001010010001110111010000110101100011101100000010010011110010011101101001111101010001011101000001011100000001100100010101110000110101110011000001001001110001101101010100011101110001100011011110001010101100000010010100101101010011100111100100110011011010000000011011110010000011001101001011011001111000010001111101011011110011011001001000000110011100011100110101110101111110111000110010011010000110100001110011110001011100011001111111000011011111011001000011111010011110100011111100100011110111010011010111110000011100011010100010111111000000010111100111001100111111001000011001000111110010000011011110011101000111000110101111100010000011101111111100000011111001011001100101101111101001100010110011101100011100101110011111011010110100001010010011011100110000001100000010111100101011011101000111101001100101101000101100101111011000000101011001000111001101100111111111111001010101100010010100101110111100111110110010100111011101010100111001000110001001000111100011111110111100100000101000000110011111110011010110111001101100000100011111011010000111100011110010111011101010110111100100000111110100100001111011101111101111001001101010010001100111000001010000010;
	localparam PROTOTYPE_A_LOW  =   2000'b10010011001110100010101101010000110100101010011001110100000101100111010101110111000001110010011100010111000111000010110010111111101000001100111111010011010010001001000000010011110010100110101010010011111101001101100001000110101111100100110011100000100011001100100100110111010011000101010011101001010111011011010111001111111000110001101000010011001111001100101100111001011000011000011100000111001010000100100111111101010100000101101101101011000001111001110111001110101111100001110111010110100000110011011001101010110001010100000101010011110110011000110001010010100111011101111010001011101110111010110000100000110101111100011001000110001110001001100011000110010100110100001011011011111100010000000110011101111110111010100011100011100011001010111100011001001011111101111011011111001000011011010010001011001000010000111101000011101100001010011001000001010010001110111010000110101100011101111100010010101110011101101101001111111110001011101000001011100000001100100010110010010110101110011000000111001110001101101010100011101110001100011011110001100101110000010010011101101010011010000100100110000111010010000011011110010000011001101001000011001111000010001111101011010000011011001001000000110001100011100110101110101111110111001000011101110000000100001110011110001011100100000011111000011011111011001000011111011100001001101111100100011110110000011010111110000011100011010100000111111000000010111100111001100111111001000100001001011110010000011011110011101000111000110101111100010000011101111111100000011111101011001100101101100001001100010110011101100011100101110011111011011000100001010010011011100110000001110000010111100101011000001000111101001100111101011101100101110001000110011011110000000010001100111110111111001010101100010010100110010110010111110110010100111011010010100111001011110000111000111100011010110111100100100100000000110011111110011011010000001101100000100011111011010000111100011110010111011101010110111101100000111110111000001111011110111101111001001101010010001100111000001010000010;
 
	hv_binary_adder #(
		.AM_NUM_FOLDS          (AM_NUM_FOLDS),
		.AM_NUM_FOLDS_WIDTH    (AM_NUM_FOLDS_WIDTH), 
		.AM_FOLD_WIDTH         (AM_FOLD_WIDTH) 
    ) BIN_ADDER (
		.hv			(similarity_hv),
		.distance	(distance)
	);

	assign hvin_fire 	= hvin_valid && hvin_ready;
	assign hvin_ready	= prototype_counter == 0 && fold_counter == 0;

	assign dout_fire 	= dout_valid && dout_ready;
	assign dout_valid	= prototype_counter == 4;
 
	always @(posedge clk) begin
		if (rst || dout_fire)
			prototype_counter <= 0;
		else if (fold_counter == AM_NUM_FOLDS-1)
			prototype_counter <= prototype_counter + 1;
	end

	always @(posedge clk) begin
		if (rst || fold_counter == AM_NUM_FOLDS-1 || dout_fire)
			fold_counter <= 0;
		else if (hvin_fire || (fold_counter > 0 && fold_counter < AM_NUM_FOLDS-1) ||
				(fold_counter == 0 && prototype_counter > 0 && prototype_counter < 4))
			fold_counter <= fold_counter + 1;
	end

	always @(*) begin
		if (prototype_counter == 0) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_V_PLUS[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
		else if (prototype_counter == 1) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_V_MIN[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
		else if (prototype_counter == 2) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_A_HIGH[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
		else if (prototype_counter == 3) begin
			similarity_hv = hvin[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH] ^ PROTOTYPE_A_LOW[(fold_counter * AM_FOLD_WIDTH) +: AM_FOLD_WIDTH];
		end
	end

	always @(posedge clk) begin
		if (prototype_counter == 0 || prototype_counter == 2) begin
			if (fold_counter == 0) 
				distance_p <= distance;
			else
				distance_p <= distance_p + distance;
		end		
	end

	always @(posedge clk) begin
		if (prototype_counter == 1 || prototype_counter == 3) begin
			if (fold_counter == 0) 
				distance_n <= distance;
			else
				distance_n <= distance_n + distance;
		end		
	end

	always @(posedge clk) begin
		if (prototype_counter == 1 && fold_counter == AM_NUM_FOLDS-1) begin
			valence <= distance_p >= (distance_n + distance);
		end

		if (prototype_counter == 3 && fold_counter == AM_NUM_FOLDS-1) begin
			arousal <= distance_p >= (distance_n + distance);
		end
	end

endmodule : associative_memory
