`ifndef CONST
`define CONST

`define HV_DIMENSION 2000
`define CHANNEL_WIDTH 2
`define NGRAM_SIZE 3
`define TOTAL_NUM_CHANNEL 214
`define GSR_SRAM_ADDR_WIDTH 5
`define ECG_SRAM_ADDR_WIDTH 7
`define EEG_SRAM_ADDR_WIDTH 7
`define GSR_NUM_CHANNEL 32
`define ECG_NUM_CHANNEL 77
`define EEG_NUM_CHANNEL 105

`define ceilLog2(x) ( \
(x) > 2**30 ? 31 : \
(x) > 2**29 ? 30 : \
(x) > 2**28 ? 29 : \
(x) > 2**27 ? 28 : \
(x) > 2**26 ? 27 : \
(x) > 2**25 ? 26 : \
(x) > 2**24 ? 25 : \
(x) > 2**23 ? 24 : \
(x) > 2**22 ? 23 : \
(x) > 2**21 ? 22 : \
(x) > 2**20 ? 21 : \
(x) > 2**19 ? 20 : \
(x) > 2**18 ? 19 : \
(x) > 2**17 ? 18 : \
(x) > 2**16 ? 17 : \
(x) > 2**15 ? 16 : \
(x) > 2**14 ? 15 : \
(x) > 2**13 ? 14 : \
(x) > 2**12 ? 13 : \
(x) > 2**11 ? 12 : \
(x) > 2**10 ? 11 : \
(x) > 2**9 ? 10 : \
(x) > 2**8 ? 9 : \
(x) > 2**7 ? 8 : \
(x) > 2**6 ? 7 : \
(x) > 2**5 ? 6 : \
(x) > 2**4 ? 5 : \
(x) > 2**3 ? 4 : \
(x) > 2**2 ? 3 : \
(x) > 2**1 ? 2 : \
(x) > 2**0 ? 1 : 0)

`define PROTOTYPE_V_PLUS 2000'b10111010111000001100110110000000111001010101110010010001111010101110100010110000111110111001010010000101000110000000001010011110000111011000101010101001011111001100110010001110100111000100011100011011011000111010111000101100000010001001000110101000001000010101101010110011100000010000000110110110100101010001010011101101111000001010000000110011110111111111000011001011000100010100011101111111011000100100001111011000101111110100111100110100001001010000101000011110011011111010010001101011001011111111101101000100001010010011100001010000110011100100001100101011101111010101111000110111111011010111100000101001000000001100010110010100100000111000000010111100001100101111101101111001111010101100111101100111111110010101110100000011100110101001010001111101111111100010100000101010110001010100101111010110000000101011111000010101000111010100111100010110111011001101111100010101101011111010010000011011111110001011100011011011000100100110101100000111000000110110110111001101000010110000010011110111011111101101101100000100111010001010000101100110100010010111001110001001001001010000100011010011111111010001101000001001001000110011111110001110101100011101000001011000001110001101011010010001100011011001011110100110111111011001010001000110101011000110011001001110000100101111101000001110111111100010011111001101110101100110011110101100001101100100010000000111100000001110010100011011111100100100001010001000100001101010111101100011000010100000100111111000110000001001010011110011110110111000101010110100010110011110000010100111001101110111000001010111111000001011000010100111001101100110100100010001111001010001110000010010111001000101000000001101101010101111010010100111110001010001010010101111110011001001101100101111010101100110000000000110101001101111011011100011000110001011010100110011111100011010101100010100111000010001110100011011101001101101001101001011011101010001101111101101010010011100011000010011110010011100101010110111111100011000110011101000111110000010101101000010000100001010011000110110

`define PROTOTYPE_V_MIN 2000'b00101010111000001110110110000000101110011011110010010000011010101110100010110000111011111001010001000001000110000000001010011110000101011000101101101010010001001100110011101110100111000100111100011000011111111010111010000000000010001000110000101000000000010101101111110011100000011001010110110110100101010001010011101101111010001000000000110010010111111111000011001011000100001000000001111111010000100100001111011001001111110100111100110100001001010000001000011110001011111010011010101011001111111111101101000100001010010011100100110000101011100100100010101010011110100001111000000001110111010111100000100001110100001100001110000000100100111100110010111100001100101111101101111000011010101100000100000111111110010101110101010001001110101001010001111101111111100010011000101010110000010100101111101110001110101011110100010101000110110100111100010110111011001101111100000101101011100110010000011011110000000101011001011011000101000110111100110111000100100110110111001101000110010000010001110111011111101101101100000101001010001010001011001110000010010111000010001001001001010000100011110100111111010001101000001000001000100011110110000010110000011101000110011000001110001101011110011001001011011001011110100110111011011001010001011001010111000001011001001110001100010111101011001110111111100010010001000101110101100110011110101100001001110111010000000111100000001110100100001011111100100100001010110000100001110110011001100010110010100000100111001000110000001001010011110111111000111010101010110100010110011110100010100111001101110111000001010111100100011100000001100111000101101010100100010001111001001101110000010010110111000101000000101101101010101111010010100110010001111011010010101111001111001000101101001100110101100111100000011010101010001100011011100011000100111011010100110011111101011010101100010100111000010001110100011011101001101101000001001011011101010011101111100011010010101100011000010111110010010010001010110010001100011000110011101000111110000010101101000010000100001010011001110011

`define PROTOTYPE_A_HIGH 2000'b00111010111000001100110110111000101100010101110010010001111010101110100010110000111110111001010101010101000110000000001010011110000111111000101101101011010101001100111000001110100111000100101100011011011111111010111000001100000010001000110000101000001000010101101101110011100110011001110110110110100101010001010011101101111000001001100000110011110111111111110010111011000100010100011111111111010000100100001111011000001111110100111100110100101001010001001000011110011111001010100010101010111011111111101101000100001010010011100100110000101011100100001010101010011111000101111000110111111011010111100100101001010000001100001110001000100010111100000010111100001100101111101101111001111010101100111100110111111110010101110100000001100110101001010001111101111111100010100000101010110000010100101111010110000110001011111000010101000101010100111100011110111011001101111100010101101011111110010000111011111110001011110101011011000101000110111100000111000101100110110111001101000101110000010011110111011111101101101100000101001010001010001011001110000010010111001110000001001001010000100011110011111111010001101000001000001000100001111110011110110000011101000110011000001110001101011110010111101011011001011110100110111001011001010001011001011111000110011001001110110100100111001011001110111111100010011111011101110101100110011110101100001100000100010000000111100000001110100100001011111100100100101010111000100001111110100101100011110010110000100111001000110000001001010011110011111100111010101010110100010110011110011010100111001101110111000001010111100100001111000010100111110101110110100100010001111001001101110000010010111001000101000001001101101010101111010010100111110001010111010010101111011111001001101101001100110101100111100000011110101010001100111011100011000110110001010100110011111100011010101100010100111000010010110100011011101001101101000101001000111101011101101111100011010010101100011000001111110010010010101010110010001100011000110011101000111110000010101101000010000100001010011001010111

`define PROTOTYPE_A_LOW 2000'b10101010111000001011110110001000111110110111110010010000011010101110100010110000111111111001010010000101000110000000001010111110000100011000101011101010011111001100110010001110100111000100111100011010111000111010111011100010000010001001000000101000001000010101101110110011100000010001000110110110100101010001010011101101111000001010000000110011110111111111100011001011010100011000011101111111011000100100001111011001111111110100111100110100010001010000111000011110000011111010011110101011001101111111101101000100001010010011100100110000110111100100001100101011101110100001111000010011110111010111100001101111101100001100011110010100100010111100110010111100001100101111001101111000011010101100010100000111111110010101110100001111100110101001010001111101111111100010100000101010110111010100101111100110000010101011110000010101000110110100111100010110111011001101111100001001101011111110010000011011111110000101011011011011000100110110111101000111000000110110110111001101000010110000010011110111011111101101101100000100111010001010000101100110000010010111010010001001001001010000100011110011111111010001101000001000001001110011011110000010101100011101000110011000001110001101011110010111010011011001011110100110111111011001011101011001001111000110011001001110000100011111101000001110111111100010010001111101110101100110011110101100001101110111010000000111100000001110010100010111111100100100001010110000100001100010111001100011110010101000100111101000101100001001010011110011111100111110101010110100010110011110100010100111001101110111000001010111111000101000000010100111000101101010100100010001111001010001110000010010110111011001000100001101101010100111010010100110010001010001010010101111000011001001101101001111010101100111010000000010101010001111011011100011000110000011111100110011111100011010101100010100111000010001110100011011111001101101001100001011001101010001101111101101010010101100011000010011110010011100101010110010101100011000110011101000111110000010101101000010000100001010011000110110

`endif